// Generator : SpinalHDL dev    git head : 008a72bc159840e8d5ca7ed6a07e1bdc5f0a9224
// Component : VexiiRiscvLitex_b3ea249d694d3e23c54ffbfd7a72a07a
// Git hash  : 63b6844fb4a8b9e88e9de55fc7b5113b30ab45d2

`timescale 1ns/1ps

module VexiiRiscvLitex_b3ea249d694d3e23c54ffbfd7a72a07a (
  input  wire          litex_reset,
  output wire          vexiis_0_cfuBus_node_cmd_valid,
  input  wire          vexiis_0_cfuBus_node_cmd_ready,
  output wire [2:0]    vexiis_0_cfuBus_node_cmd_payload_function_id,
  output wire [31:0]   vexiis_0_cfuBus_node_cmd_payload_inputs_0,
  output wire [31:0]   vexiis_0_cfuBus_node_cmd_payload_inputs_1,
  input  wire          vexiis_0_cfuBus_node_rsp_valid,
  output wire          vexiis_0_cfuBus_node_rsp_ready,
  input  wire [31:0]   vexiis_0_cfuBus_node_rsp_payload_outputs_0,
  input  wire [31:0]   peripheral_externalInterrupts_port,
  output wire          mBus_awvalid,
  input  wire          mBus_awready,
  output wire [31:0]   mBus_awaddr,
  output wire [7:0]    mBus_awid,
  output wire [7:0]    mBus_awlen,
  output wire [2:0]    mBus_awsize,
  output wire [1:0]    mBus_awburst,
  output wire          mBus_awallStrb,
  output wire          mBus_wvalid,
  input  wire          mBus_wready,
  output wire [127:0]  mBus_wdata,
  output wire [15:0]   mBus_wstrb,
  output wire          mBus_wlast,
  input  wire          mBus_bvalid,
  output wire          mBus_bready,
  input  wire [7:0]    mBus_bid,
  input  wire [1:0]    mBus_bresp,
  output wire          mBus_arvalid,
  input  wire          mBus_arready,
  output wire [31:0]   mBus_araddr,
  output wire [7:0]    mBus_arid,
  output wire [7:0]    mBus_arlen,
  output wire [2:0]    mBus_arsize,
  output wire [1:0]    mBus_arburst,
  input  wire          mBus_rvalid,
  output wire          mBus_rready,
  input  wire [127:0]  mBus_rdata,
  input  wire [7:0]    mBus_rid,
  input  wire [1:0]    mBus_rresp,
  input  wire          mBus_rlast,
  output wire          pBus_awvalid,
  input  wire          pBus_awready,
  output wire [31:0]   pBus_awaddr,
  output wire [2:0]    pBus_awprot,
  output wire          pBus_wvalid,
  input  wire          pBus_wready,
  output wire [31:0]   pBus_wdata,
  output wire [3:0]    pBus_wstrb,
  input  wire          pBus_bvalid,
  output wire          pBus_bready,
  input  wire [1:0]    pBus_bresp,
  output wire          pBus_arvalid,
  input  wire          pBus_arready,
  output wire [31:0]   pBus_araddr,
  output wire [2:0]    pBus_arprot,
  input  wire          pBus_rvalid,
  output wire          pBus_rready,
  input  wire [31:0]   pBus_rdata,
  input  wire [1:0]    pBus_rresp,
  output reg  [7:0]    debug,
  input  wire          litex_clk
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                peripheral_clint_thread_core_io_stop;
  reg        [30:0]   peripheral_plic_thread_logic_io_sources;
  wire                peripheral_bus_decoder_core_io_up_d_ready;
  wire                vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_valid;
  wire       [2:0]    vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_function_id;
  wire       [31:0]   vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_inputs_0;
  wire       [31:0]   vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_inputs_1;
  wire       [2:0]    vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_state_index;
  wire       [3:0]    vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_cfu_index;
  wire       [31:0]   vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_raw_insn;
  wire                vexiis_0_logic_core_CfuPlugin_logic_bus_rsp_ready;
  wire                vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_valid;
  wire       [2:0]    vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_opcode;
  wire       [2:0]    vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_param;
  wire       [31:0]   vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_address;
  wire       [2:0]    vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_size;
  wire                vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_d_ready;
  wire                vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_valid;
  wire       [2:0]    vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_opcode;
  wire       [2:0]    vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_param;
  wire       [0:0]    vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_source;
  wire       [31:0]   vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_address;
  wire       [2:0]    vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_size;
  wire       [7:0]    vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_mask;
  wire       [63:0]   vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_data;
  wire                vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_corrupt;
  wire                vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_d_ready;
  wire                vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_valid;
  wire       [2:0]    vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode;
  wire       [2:0]    vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_param;
  wire       [31:0]   vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_address;
  wire       [1:0]    vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_size;
  wire       [3:0]    vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_mask;
  wire       [31:0]   vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_data;
  wire                vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt;
  wire                vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_d_ready;
  wire                cpuResetCtrl_fiber_aggregator_asyncBuffers_0_io_dataOut;
  wire                cpuResetCtrl_fiber_buffer_io_dataOut;
  wire                splited_mBus_arbiter_core_io_ups_0_a_ready;
  wire                splited_mBus_arbiter_core_io_ups_0_d_valid;
  wire       [2:0]    splited_mBus_arbiter_core_io_ups_0_d_payload_opcode;
  wire       [2:0]    splited_mBus_arbiter_core_io_ups_0_d_payload_param;
  wire       [2:0]    splited_mBus_arbiter_core_io_ups_0_d_payload_size;
  wire                splited_mBus_arbiter_core_io_ups_0_d_payload_denied;
  wire       [63:0]   splited_mBus_arbiter_core_io_ups_0_d_payload_data;
  wire                splited_mBus_arbiter_core_io_ups_0_d_payload_corrupt;
  wire                splited_mBus_arbiter_core_io_ups_1_a_ready;
  wire                splited_mBus_arbiter_core_io_ups_1_d_valid;
  wire       [2:0]    splited_mBus_arbiter_core_io_ups_1_d_payload_opcode;
  wire       [2:0]    splited_mBus_arbiter_core_io_ups_1_d_payload_param;
  wire       [0:0]    splited_mBus_arbiter_core_io_ups_1_d_payload_source;
  wire       [2:0]    splited_mBus_arbiter_core_io_ups_1_d_payload_size;
  wire                splited_mBus_arbiter_core_io_ups_1_d_payload_denied;
  wire       [63:0]   splited_mBus_arbiter_core_io_ups_1_d_payload_data;
  wire                splited_mBus_arbiter_core_io_ups_1_d_payload_corrupt;
  wire                splited_mBus_arbiter_core_io_down_a_valid;
  wire       [2:0]    splited_mBus_arbiter_core_io_down_a_payload_opcode;
  wire       [2:0]    splited_mBus_arbiter_core_io_down_a_payload_param;
  wire       [1:0]    splited_mBus_arbiter_core_io_down_a_payload_source;
  wire       [31:0]   splited_mBus_arbiter_core_io_down_a_payload_address;
  wire       [2:0]    splited_mBus_arbiter_core_io_down_a_payload_size;
  wire       [7:0]    splited_mBus_arbiter_core_io_down_a_payload_mask;
  wire       [63:0]   splited_mBus_arbiter_core_io_down_a_payload_data;
  wire                splited_mBus_arbiter_core_io_down_a_payload_corrupt;
  wire                splited_mBus_arbiter_core_io_down_d_ready;
  wire                peripheral_bus_arbiter_core_io_ups_0_a_ready;
  wire                peripheral_bus_arbiter_core_io_ups_0_d_valid;
  wire       [2:0]    peripheral_bus_arbiter_core_io_ups_0_d_payload_opcode;
  wire       [2:0]    peripheral_bus_arbiter_core_io_ups_0_d_payload_param;
  wire       [1:0]    peripheral_bus_arbiter_core_io_ups_0_d_payload_size;
  wire                peripheral_bus_arbiter_core_io_ups_0_d_payload_denied;
  wire       [31:0]   peripheral_bus_arbiter_core_io_ups_0_d_payload_data;
  wire                peripheral_bus_arbiter_core_io_ups_0_d_payload_corrupt;
  wire                peripheral_bus_arbiter_core_io_ups_1_a_ready;
  wire                peripheral_bus_arbiter_core_io_ups_1_d_valid;
  wire       [2:0]    peripheral_bus_arbiter_core_io_ups_1_d_payload_opcode;
  wire       [2:0]    peripheral_bus_arbiter_core_io_ups_1_d_payload_param;
  wire       [1:0]    peripheral_bus_arbiter_core_io_ups_1_d_payload_source;
  wire       [2:0]    peripheral_bus_arbiter_core_io_ups_1_d_payload_size;
  wire                peripheral_bus_arbiter_core_io_ups_1_d_payload_denied;
  wire       [31:0]   peripheral_bus_arbiter_core_io_ups_1_d_payload_data;
  wire                peripheral_bus_arbiter_core_io_ups_1_d_payload_corrupt;
  wire                peripheral_bus_arbiter_core_io_down_a_valid;
  wire       [2:0]    peripheral_bus_arbiter_core_io_down_a_payload_opcode;
  wire       [2:0]    peripheral_bus_arbiter_core_io_down_a_payload_param;
  wire       [2:0]    peripheral_bus_arbiter_core_io_down_a_payload_source;
  wire       [31:0]   peripheral_bus_arbiter_core_io_down_a_payload_address;
  wire       [2:0]    peripheral_bus_arbiter_core_io_down_a_payload_size;
  wire       [3:0]    peripheral_bus_arbiter_core_io_down_a_payload_mask;
  wire       [31:0]   peripheral_bus_arbiter_core_io_down_a_payload_data;
  wire                peripheral_bus_arbiter_core_io_down_a_payload_corrupt;
  wire                peripheral_bus_arbiter_core_io_down_d_ready;
  wire                mem_toAxi4_logic_bridge_io_up_a_ready;
  wire                mem_toAxi4_logic_bridge_io_up_d_valid;
  wire       [2:0]    mem_toAxi4_logic_bridge_io_up_d_payload_opcode;
  wire       [2:0]    mem_toAxi4_logic_bridge_io_up_d_payload_param;
  wire       [1:0]    mem_toAxi4_logic_bridge_io_up_d_payload_source;
  wire       [2:0]    mem_toAxi4_logic_bridge_io_up_d_payload_size;
  wire                mem_toAxi4_logic_bridge_io_up_d_payload_denied;
  wire       [127:0]  mem_toAxi4_logic_bridge_io_up_d_payload_data;
  wire                mem_toAxi4_logic_bridge_io_up_d_payload_corrupt;
  wire                mem_toAxi4_logic_bridge_io_down_ar_valid;
  wire       [31:0]   mem_toAxi4_logic_bridge_io_down_ar_payload_addr;
  wire       [1:0]    mem_toAxi4_logic_bridge_io_down_ar_payload_id;
  wire       [7:0]    mem_toAxi4_logic_bridge_io_down_ar_payload_len;
  wire       [2:0]    mem_toAxi4_logic_bridge_io_down_ar_payload_size;
  wire       [1:0]    mem_toAxi4_logic_bridge_io_down_ar_payload_burst;
  wire                mem_toAxi4_logic_bridge_io_down_aw_valid;
  wire       [31:0]   mem_toAxi4_logic_bridge_io_down_aw_payload_addr;
  wire       [1:0]    mem_toAxi4_logic_bridge_io_down_aw_payload_id;
  wire       [7:0]    mem_toAxi4_logic_bridge_io_down_aw_payload_len;
  wire       [2:0]    mem_toAxi4_logic_bridge_io_down_aw_payload_size;
  wire       [1:0]    mem_toAxi4_logic_bridge_io_down_aw_payload_burst;
  wire                mem_toAxi4_logic_bridge_io_down_aw_payload_allStrb;
  wire                mem_toAxi4_logic_bridge_io_down_w_valid;
  wire       [127:0]  mem_toAxi4_logic_bridge_io_down_w_payload_data;
  wire       [15:0]   mem_toAxi4_logic_bridge_io_down_w_payload_strb;
  wire                mem_toAxi4_logic_bridge_io_down_w_payload_last;
  wire                mem_toAxi4_logic_bridge_io_down_r_ready;
  wire                mem_toAxi4_logic_bridge_io_down_b_ready;
  wire                splited_mBus_decoder_core_io_up_a_ready;
  wire                splited_mBus_decoder_core_io_up_d_valid;
  wire       [2:0]    splited_mBus_decoder_core_io_up_d_payload_opcode;
  wire       [2:0]    splited_mBus_decoder_core_io_up_d_payload_param;
  wire       [1:0]    splited_mBus_decoder_core_io_up_d_payload_source;
  wire       [2:0]    splited_mBus_decoder_core_io_up_d_payload_size;
  wire                splited_mBus_decoder_core_io_up_d_payload_denied;
  wire       [63:0]   splited_mBus_decoder_core_io_up_d_payload_data;
  wire                splited_mBus_decoder_core_io_up_d_payload_corrupt;
  wire                splited_mBus_decoder_core_io_downs_0_a_valid;
  wire       [2:0]    splited_mBus_decoder_core_io_downs_0_a_payload_opcode;
  wire       [2:0]    splited_mBus_decoder_core_io_downs_0_a_payload_param;
  wire       [1:0]    splited_mBus_decoder_core_io_downs_0_a_payload_source;
  wire       [31:0]   splited_mBus_decoder_core_io_downs_0_a_payload_address;
  wire       [2:0]    splited_mBus_decoder_core_io_downs_0_a_payload_size;
  wire       [7:0]    splited_mBus_decoder_core_io_downs_0_a_payload_mask;
  wire       [63:0]   splited_mBus_decoder_core_io_downs_0_a_payload_data;
  wire                splited_mBus_decoder_core_io_downs_0_a_payload_corrupt;
  wire                splited_mBus_decoder_core_io_downs_0_d_ready;
  wire                splited_mBus_decoder_core_io_downs_1_a_valid;
  wire       [2:0]    splited_mBus_decoder_core_io_downs_1_a_payload_opcode;
  wire       [2:0]    splited_mBus_decoder_core_io_downs_1_a_payload_param;
  wire       [1:0]    splited_mBus_decoder_core_io_downs_1_a_payload_source;
  wire       [31:0]   splited_mBus_decoder_core_io_downs_1_a_payload_address;
  wire       [2:0]    splited_mBus_decoder_core_io_downs_1_a_payload_size;
  wire       [7:0]    splited_mBus_decoder_core_io_downs_1_a_payload_mask;
  wire       [63:0]   splited_mBus_decoder_core_io_downs_1_a_payload_data;
  wire                splited_mBus_decoder_core_io_downs_1_a_payload_corrupt;
  wire                splited_mBus_decoder_core_io_downs_1_d_ready;
  wire                peripheral_clint_thread_core_io_bus_a_ready;
  wire                peripheral_clint_thread_core_io_bus_d_valid;
  wire       [2:0]    peripheral_clint_thread_core_io_bus_d_payload_opcode;
  wire       [2:0]    peripheral_clint_thread_core_io_bus_d_payload_param;
  wire       [2:0]    peripheral_clint_thread_core_io_bus_d_payload_source;
  wire       [2:0]    peripheral_clint_thread_core_io_bus_d_payload_size;
  wire                peripheral_clint_thread_core_io_bus_d_payload_denied;
  wire       [31:0]   peripheral_clint_thread_core_io_bus_d_payload_data;
  wire                peripheral_clint_thread_core_io_bus_d_payload_corrupt;
  wire       [0:0]    peripheral_clint_thread_core_io_timerInterrupt;
  wire       [0:0]    peripheral_clint_thread_core_io_softwareInterrupt;
  wire       [63:0]   peripheral_clint_thread_core_io_time;
  wire                peripheral_plic_thread_logic_io_bus_a_ready;
  wire                peripheral_plic_thread_logic_io_bus_d_valid;
  wire       [2:0]    peripheral_plic_thread_logic_io_bus_d_payload_opcode;
  wire       [2:0]    peripheral_plic_thread_logic_io_bus_d_payload_param;
  wire       [2:0]    peripheral_plic_thread_logic_io_bus_d_payload_source;
  wire       [1:0]    peripheral_plic_thread_logic_io_bus_d_payload_size;
  wire                peripheral_plic_thread_logic_io_bus_d_payload_denied;
  wire       [31:0]   peripheral_plic_thread_logic_io_bus_d_payload_data;
  wire                peripheral_plic_thread_logic_io_bus_d_payload_corrupt;
  wire       [1:0]    peripheral_plic_thread_logic_io_targets;
  wire                peripheral_toAxiLite4_logic_bridge_io_up_a_ready;
  wire                peripheral_toAxiLite4_logic_bridge_io_up_d_valid;
  wire       [2:0]    peripheral_toAxiLite4_logic_bridge_io_up_d_payload_opcode;
  wire       [2:0]    peripheral_toAxiLite4_logic_bridge_io_up_d_payload_param;
  wire       [2:0]    peripheral_toAxiLite4_logic_bridge_io_up_d_payload_source;
  wire       [2:0]    peripheral_toAxiLite4_logic_bridge_io_up_d_payload_size;
  wire                peripheral_toAxiLite4_logic_bridge_io_up_d_payload_denied;
  wire       [31:0]   peripheral_toAxiLite4_logic_bridge_io_up_d_payload_data;
  wire                peripheral_toAxiLite4_logic_bridge_io_up_d_payload_corrupt;
  wire                peripheral_toAxiLite4_logic_bridge_io_down_aw_valid;
  wire       [31:0]   peripheral_toAxiLite4_logic_bridge_io_down_aw_payload_addr;
  wire       [2:0]    peripheral_toAxiLite4_logic_bridge_io_down_aw_payload_prot;
  wire                peripheral_toAxiLite4_logic_bridge_io_down_w_valid;
  wire       [31:0]   peripheral_toAxiLite4_logic_bridge_io_down_w_payload_data;
  wire       [3:0]    peripheral_toAxiLite4_logic_bridge_io_down_w_payload_strb;
  wire                peripheral_toAxiLite4_logic_bridge_io_down_b_ready;
  wire                peripheral_toAxiLite4_logic_bridge_io_down_ar_valid;
  wire       [31:0]   peripheral_toAxiLite4_logic_bridge_io_down_ar_payload_addr;
  wire       [2:0]    peripheral_toAxiLite4_logic_bridge_io_down_ar_payload_prot;
  wire                peripheral_toAxiLite4_logic_bridge_io_down_r_ready;
  wire                splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_a_ready;
  wire                splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_valid;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_opcode;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_param;
  wire       [1:0]    splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_source;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_size;
  wire                splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_denied;
  wire       [63:0]   splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_data;
  wire                splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_corrupt;
  wire                splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_valid;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_opcode;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_param;
  wire       [1:0]    splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_source;
  wire       [31:0]   splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_address;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_size;
  wire       [15:0]   splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_mask;
  wire       [127:0]  splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_data;
  wire                splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_corrupt;
  wire                splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_d_ready;
  wire                splited_mBus_to_peripheral_bus_widthAdapter_io_up_a_ready;
  wire                splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_valid;
  wire       [2:0]    splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_opcode;
  wire       [2:0]    splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_param;
  wire       [1:0]    splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_source;
  wire       [2:0]    splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_size;
  wire                splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_denied;
  wire       [63:0]   splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_data;
  wire                splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_corrupt;
  wire                splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_valid;
  wire       [2:0]    splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_opcode;
  wire       [2:0]    splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_param;
  wire       [1:0]    splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_source;
  wire       [31:0]   splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_address;
  wire       [2:0]    splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_size;
  wire       [3:0]    splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_mask;
  wire       [31:0]   splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_data;
  wire                splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_corrupt;
  wire                splited_mBus_to_peripheral_bus_widthAdapter_io_down_d_ready;
  wire                peripheral_bus_decoder_core_io_up_a_ready;
  wire                peripheral_bus_decoder_core_io_up_d_valid;
  wire       [2:0]    peripheral_bus_decoder_core_io_up_d_payload_opcode;
  wire       [2:0]    peripheral_bus_decoder_core_io_up_d_payload_param;
  wire       [2:0]    peripheral_bus_decoder_core_io_up_d_payload_source;
  wire       [2:0]    peripheral_bus_decoder_core_io_up_d_payload_size;
  wire                peripheral_bus_decoder_core_io_up_d_payload_denied;
  wire       [31:0]   peripheral_bus_decoder_core_io_up_d_payload_data;
  wire                peripheral_bus_decoder_core_io_up_d_payload_corrupt;
  wire                peripheral_bus_decoder_core_io_downs_0_a_valid;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_0_a_payload_opcode;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_0_a_payload_param;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_0_a_payload_source;
  wire       [15:0]   peripheral_bus_decoder_core_io_downs_0_a_payload_address;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_0_a_payload_size;
  wire       [3:0]    peripheral_bus_decoder_core_io_downs_0_a_payload_mask;
  wire       [31:0]   peripheral_bus_decoder_core_io_downs_0_a_payload_data;
  wire                peripheral_bus_decoder_core_io_downs_0_a_payload_corrupt;
  wire                peripheral_bus_decoder_core_io_downs_0_d_ready;
  wire                peripheral_bus_decoder_core_io_downs_1_a_valid;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_1_a_payload_opcode;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_1_a_payload_param;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_1_a_payload_source;
  wire       [21:0]   peripheral_bus_decoder_core_io_downs_1_a_payload_address;
  wire       [1:0]    peripheral_bus_decoder_core_io_downs_1_a_payload_size;
  wire       [3:0]    peripheral_bus_decoder_core_io_downs_1_a_payload_mask;
  wire       [31:0]   peripheral_bus_decoder_core_io_downs_1_a_payload_data;
  wire                peripheral_bus_decoder_core_io_downs_1_a_payload_corrupt;
  wire                peripheral_bus_decoder_core_io_downs_1_d_ready;
  wire                peripheral_bus_decoder_core_io_downs_2_a_valid;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_2_a_payload_opcode;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_2_a_payload_param;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_2_a_payload_source;
  wire       [31:0]   peripheral_bus_decoder_core_io_downs_2_a_payload_address;
  wire       [2:0]    peripheral_bus_decoder_core_io_downs_2_a_payload_size;
  wire       [3:0]    peripheral_bus_decoder_core_io_downs_2_a_payload_mask;
  wire       [31:0]   peripheral_bus_decoder_core_io_downs_2_a_payload_data;
  wire                peripheral_bus_decoder_core_io_downs_2_a_payload_corrupt;
  wire                peripheral_bus_decoder_core_io_downs_2_d_ready;
  wire                cpuResetCtrl_reset;
  wire       [2:0]    vexiis_0_cfuBus_node_cmd_payload_state_index;
  wire       [3:0]    vexiis_0_cfuBus_node_cmd_payload_cfu_index;
  wire       [31:0]   vexiis_0_cfuBus_node_cmd_payload_raw_insn;
  wire                vexiis_0_priv_mti_flag;
  wire                vexiis_0_priv_msi_flag;
  wire                vexiis_0_priv_mei_flag;
  wire                vexiis_0_priv_sei_flag;
  wire                vexiis_0_priv_stoptime;
  wire       [63:0]   vexiis_0_priv_rdtime;
  wire       [63:0]   peripheral_clint_time;
  wire                peripheral_externalInterrupts_toPlic_1_node_flag;
  wire                peripheral_externalInterrupts_toPlic_2_node_flag;
  wire                peripheral_externalInterrupts_toPlic_3_node_flag;
  wire                peripheral_externalInterrupts_toPlic_4_node_flag;
  wire                peripheral_externalInterrupts_toPlic_5_node_flag;
  wire                peripheral_externalInterrupts_toPlic_6_node_flag;
  wire                peripheral_externalInterrupts_toPlic_7_node_flag;
  wire                peripheral_externalInterrupts_toPlic_8_node_flag;
  wire                peripheral_externalInterrupts_toPlic_9_node_flag;
  wire                peripheral_externalInterrupts_toPlic_10_node_flag;
  wire                peripheral_externalInterrupts_toPlic_11_node_flag;
  wire                peripheral_externalInterrupts_toPlic_12_node_flag;
  wire                peripheral_externalInterrupts_toPlic_13_node_flag;
  wire                peripheral_externalInterrupts_toPlic_14_node_flag;
  wire                peripheral_externalInterrupts_toPlic_15_node_flag;
  wire                peripheral_externalInterrupts_toPlic_16_node_flag;
  wire                peripheral_externalInterrupts_toPlic_17_node_flag;
  wire                peripheral_externalInterrupts_toPlic_18_node_flag;
  wire                peripheral_externalInterrupts_toPlic_19_node_flag;
  wire                peripheral_externalInterrupts_toPlic_20_node_flag;
  wire                peripheral_externalInterrupts_toPlic_21_node_flag;
  wire                peripheral_externalInterrupts_toPlic_22_node_flag;
  wire                peripheral_externalInterrupts_toPlic_23_node_flag;
  wire                peripheral_externalInterrupts_toPlic_24_node_flag;
  wire                peripheral_externalInterrupts_toPlic_25_node_flag;
  wire                peripheral_externalInterrupts_toPlic_26_node_flag;
  wire                peripheral_externalInterrupts_toPlic_27_node_flag;
  wire                peripheral_externalInterrupts_toPlic_28_node_flag;
  wire                peripheral_externalInterrupts_toPlic_29_node_flag;
  wire                peripheral_externalInterrupts_toPlic_30_node_flag;
  wire                peripheral_externalInterrupts_toPlic_31_node_flag;
  reg                 vexiis_0_priv_stoptime_regNext;
  reg        [63:0]   _zz_vexiis_0_priv_rdtime;
  wire                peripheral_plic_to_vexiis_0_priv_mei_flag;
  wire                peripheral_plic_to_vexiis_0_priv_sei_flag;
  wire                cpuResetCtrl_fiber_aggregator_reset;
  reg        [6:0]    cpuResetCtrl_fiber_holder_counter;
  wire                cpuResetCtrl_fiber_holder_reset;
  wire                when_CrossClock_l341;
  wire                vexiis_0_priv_mti_thread_gateways_0_flag;
  wire                vexiis_0_priv_msi_thread_gateways_0_flag;
  wire                vexiis_0_priv_mei_thread_gateways_0_flag;
  wire                vexiis_0_priv_sei_thread_gateways_0_flag;
  wire                vexiis_0_dBus_bus_a_valid;
  wire                vexiis_0_dBus_bus_a_ready;
  wire       [2:0]    vexiis_0_dBus_bus_a_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_bus_a_payload_param;
  wire       [31:0]   vexiis_0_dBus_bus_a_payload_address;
  wire       [1:0]    vexiis_0_dBus_bus_a_payload_size;
  wire       [3:0]    vexiis_0_dBus_bus_a_payload_mask;
  wire       [31:0]   vexiis_0_dBus_bus_a_payload_data;
  wire                vexiis_0_dBus_bus_a_payload_corrupt;
  wire                vexiis_0_dBus_bus_d_valid;
  wire                vexiis_0_dBus_bus_d_ready;
  wire       [2:0]    vexiis_0_dBus_bus_d_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_bus_d_payload_param;
  wire       [1:0]    vexiis_0_dBus_bus_d_payload_size;
  wire                vexiis_0_dBus_bus_d_payload_denied;
  wire       [31:0]   vexiis_0_dBus_bus_d_payload_data;
  wire                vexiis_0_dBus_bus_d_payload_corrupt;
  wire                vexiis_0_dBus_noDecoder_toDown_a_valid;
  wire                vexiis_0_dBus_noDecoder_toDown_a_ready;
  wire       [2:0]    vexiis_0_dBus_noDecoder_toDown_a_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_noDecoder_toDown_a_payload_param;
  wire       [31:0]   vexiis_0_dBus_noDecoder_toDown_a_payload_address;
  wire       [1:0]    vexiis_0_dBus_noDecoder_toDown_a_payload_size;
  wire       [3:0]    vexiis_0_dBus_noDecoder_toDown_a_payload_mask;
  wire       [31:0]   vexiis_0_dBus_noDecoder_toDown_a_payload_data;
  wire                vexiis_0_dBus_noDecoder_toDown_a_payload_corrupt;
  wire                vexiis_0_dBus_noDecoder_toDown_d_valid;
  reg                 vexiis_0_dBus_noDecoder_toDown_d_ready;
  wire       [2:0]    vexiis_0_dBus_noDecoder_toDown_d_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_noDecoder_toDown_d_payload_param;
  wire       [1:0]    vexiis_0_dBus_noDecoder_toDown_d_payload_size;
  wire                vexiis_0_dBus_noDecoder_toDown_d_payload_denied;
  wire       [31:0]   vexiis_0_dBus_noDecoder_toDown_d_payload_data;
  wire                vexiis_0_dBus_noDecoder_toDown_d_payload_corrupt;
  wire                vexiis_0_dBus_bus_a_halfPipe_valid;
  wire                vexiis_0_dBus_bus_a_halfPipe_ready;
  wire       [2:0]    vexiis_0_dBus_bus_a_halfPipe_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_bus_a_halfPipe_payload_param;
  wire       [31:0]   vexiis_0_dBus_bus_a_halfPipe_payload_address;
  wire       [1:0]    vexiis_0_dBus_bus_a_halfPipe_payload_size;
  wire       [3:0]    vexiis_0_dBus_bus_a_halfPipe_payload_mask;
  wire       [31:0]   vexiis_0_dBus_bus_a_halfPipe_payload_data;
  wire                vexiis_0_dBus_bus_a_halfPipe_payload_corrupt;
  reg                 vexiis_0_dBus_bus_a_rValid;
  wire                vexiis_0_dBus_bus_a_halfPipe_fire;
  reg        [2:0]    vexiis_0_dBus_bus_a_rData_opcode;
  reg        [2:0]    vexiis_0_dBus_bus_a_rData_param;
  reg        [31:0]   vexiis_0_dBus_bus_a_rData_address;
  reg        [1:0]    vexiis_0_dBus_bus_a_rData_size;
  reg        [3:0]    vexiis_0_dBus_bus_a_rData_mask;
  reg        [31:0]   vexiis_0_dBus_bus_a_rData_data;
  reg                 vexiis_0_dBus_bus_a_rData_corrupt;
  wire                vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_valid;
  wire                vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_ready;
  wire       [2:0]    vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_param;
  wire       [1:0]    vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_size;
  wire                vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_denied;
  wire       [31:0]   vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_data;
  wire                vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_corrupt;
  (* keep , syn_keep *) reg                 vexiis_0_dBus_noDecoder_toDown_d_rValid /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    vexiis_0_dBus_noDecoder_toDown_d_rData_opcode /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    vexiis_0_dBus_noDecoder_toDown_d_rData_param /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [1:0]    vexiis_0_dBus_noDecoder_toDown_d_rData_size /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg                 vexiis_0_dBus_noDecoder_toDown_d_rData_denied /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   vexiis_0_dBus_noDecoder_toDown_d_rData_data /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg                 vexiis_0_dBus_noDecoder_toDown_d_rData_corrupt /* synthesis syn_keep = 1 */ ;
  wire                when_Stream_l399;
  wire                vexiis_0_iBus_bus_a_valid;
  wire                vexiis_0_iBus_bus_a_ready;
  wire       [2:0]    vexiis_0_iBus_bus_a_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_bus_a_payload_param;
  wire       [31:0]   vexiis_0_iBus_bus_a_payload_address;
  wire       [2:0]    vexiis_0_iBus_bus_a_payload_size;
  wire                vexiis_0_iBus_bus_d_valid;
  wire                vexiis_0_iBus_bus_d_ready;
  wire       [2:0]    vexiis_0_iBus_bus_d_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_bus_d_payload_param;
  wire       [2:0]    vexiis_0_iBus_bus_d_payload_size;
  wire                vexiis_0_iBus_bus_d_payload_denied;
  wire       [63:0]   vexiis_0_iBus_bus_d_payload_data;
  wire                vexiis_0_iBus_bus_d_payload_corrupt;
  wire                vexiis_0_iBus_noDecoder_toDown_a_valid;
  wire                vexiis_0_iBus_noDecoder_toDown_a_ready;
  wire       [2:0]    vexiis_0_iBus_noDecoder_toDown_a_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_noDecoder_toDown_a_payload_param;
  wire       [31:0]   vexiis_0_iBus_noDecoder_toDown_a_payload_address;
  wire       [2:0]    vexiis_0_iBus_noDecoder_toDown_a_payload_size;
  wire                vexiis_0_iBus_noDecoder_toDown_d_valid;
  reg                 vexiis_0_iBus_noDecoder_toDown_d_ready;
  wire       [2:0]    vexiis_0_iBus_noDecoder_toDown_d_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_noDecoder_toDown_d_payload_param;
  wire       [2:0]    vexiis_0_iBus_noDecoder_toDown_d_payload_size;
  wire                vexiis_0_iBus_noDecoder_toDown_d_payload_denied;
  wire       [63:0]   vexiis_0_iBus_noDecoder_toDown_d_payload_data;
  wire                vexiis_0_iBus_noDecoder_toDown_d_payload_corrupt;
  wire                vexiis_0_iBus_bus_a_halfPipe_valid;
  wire                vexiis_0_iBus_bus_a_halfPipe_ready;
  wire       [2:0]    vexiis_0_iBus_bus_a_halfPipe_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_bus_a_halfPipe_payload_param;
  wire       [31:0]   vexiis_0_iBus_bus_a_halfPipe_payload_address;
  wire       [2:0]    vexiis_0_iBus_bus_a_halfPipe_payload_size;
  reg                 vexiis_0_iBus_bus_a_rValid;
  wire                vexiis_0_iBus_bus_a_halfPipe_fire;
  reg        [2:0]    vexiis_0_iBus_bus_a_rData_opcode;
  reg        [2:0]    vexiis_0_iBus_bus_a_rData_param;
  reg        [31:0]   vexiis_0_iBus_bus_a_rData_address;
  reg        [2:0]    vexiis_0_iBus_bus_a_rData_size;
  wire                vexiis_0_iBus_bus_a_halfPipe_halfPipe_valid;
  wire                vexiis_0_iBus_bus_a_halfPipe_halfPipe_ready;
  wire       [2:0]    vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_param;
  wire       [31:0]   vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_address;
  wire       [2:0]    vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_size;
  reg                 vexiis_0_iBus_bus_a_halfPipe_rValid;
  wire                vexiis_0_iBus_bus_a_halfPipe_halfPipe_fire;
  reg        [2:0]    vexiis_0_iBus_bus_a_halfPipe_rData_opcode;
  reg        [2:0]    vexiis_0_iBus_bus_a_halfPipe_rData_param;
  reg        [31:0]   vexiis_0_iBus_bus_a_halfPipe_rData_address;
  reg        [2:0]    vexiis_0_iBus_bus_a_halfPipe_rData_size;
  wire                vexiis_0_iBus_noDecoder_connection_valid;
  wire                vexiis_0_iBus_noDecoder_connection_ready;
  wire       [2:0]    vexiis_0_iBus_noDecoder_connection_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_noDecoder_connection_payload_param;
  wire       [2:0]    vexiis_0_iBus_noDecoder_connection_payload_size;
  wire                vexiis_0_iBus_noDecoder_connection_payload_denied;
  wire       [63:0]   vexiis_0_iBus_noDecoder_connection_payload_data;
  wire                vexiis_0_iBus_noDecoder_connection_payload_corrupt;
  reg                 vexiis_0_iBus_noDecoder_toDown_d_rValid;
  reg        [2:0]    vexiis_0_iBus_noDecoder_toDown_d_rData_opcode;
  reg        [2:0]    vexiis_0_iBus_noDecoder_toDown_d_rData_param;
  reg        [2:0]    vexiis_0_iBus_noDecoder_toDown_d_rData_size;
  reg                 vexiis_0_iBus_noDecoder_toDown_d_rData_denied;
  reg        [63:0]   vexiis_0_iBus_noDecoder_toDown_d_rData_data;
  reg                 vexiis_0_iBus_noDecoder_toDown_d_rData_corrupt;
  wire                when_Stream_l399_1;
  wire                vexiis_0_lsuL1Bus_bus_a_valid;
  wire                vexiis_0_lsuL1Bus_bus_a_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_a_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_a_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_bus_a_payload_source;
  wire       [31:0]   vexiis_0_lsuL1Bus_bus_a_payload_address;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_a_payload_size;
  wire       [7:0]    vexiis_0_lsuL1Bus_bus_a_payload_mask;
  wire       [63:0]   vexiis_0_lsuL1Bus_bus_a_payload_data;
  wire                vexiis_0_lsuL1Bus_bus_a_payload_corrupt;
  wire                vexiis_0_lsuL1Bus_bus_d_valid;
  wire                vexiis_0_lsuL1Bus_bus_d_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_d_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_d_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_bus_d_payload_source;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_d_payload_size;
  wire                vexiis_0_lsuL1Bus_bus_d_payload_denied;
  wire       [63:0]   vexiis_0_lsuL1Bus_bus_d_payload_data;
  wire                vexiis_0_lsuL1Bus_bus_d_payload_corrupt;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_a_valid;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_a_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_source;
  wire       [31:0]   vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_address;
  wire       [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_size;
  wire       [7:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_mask;
  wire       [63:0]   vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_data;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_corrupt;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_d_valid;
  reg                 vexiis_0_lsuL1Bus_noDecoder_toDown_d_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_source;
  wire       [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_size;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_denied;
  wire       [63:0]   vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_data;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_corrupt;
  wire                vexiis_0_lsuL1Bus_bus_a_s2mPipe_valid;
  reg                 vexiis_0_lsuL1Bus_bus_a_s2mPipe_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_source;
  wire       [31:0]   vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_address;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_size;
  wire       [7:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_mask;
  wire       [63:0]   vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_data;
  wire                vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_corrupt;
  reg                 vexiis_0_lsuL1Bus_bus_a_rValidN;
  reg        [2:0]    vexiis_0_lsuL1Bus_bus_a_rData_opcode;
  reg        [2:0]    vexiis_0_lsuL1Bus_bus_a_rData_param;
  reg        [0:0]    vexiis_0_lsuL1Bus_bus_a_rData_source;
  reg        [31:0]   vexiis_0_lsuL1Bus_bus_a_rData_address;
  reg        [2:0]    vexiis_0_lsuL1Bus_bus_a_rData_size;
  reg        [7:0]    vexiis_0_lsuL1Bus_bus_a_rData_mask;
  reg        [63:0]   vexiis_0_lsuL1Bus_bus_a_rData_data;
  reg                 vexiis_0_lsuL1Bus_bus_a_rData_corrupt;
  wire       [2:0]    _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode;
  wire                vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_valid;
  wire                vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_source;
  wire       [31:0]   vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_address;
  wire       [2:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_size;
  wire       [7:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_mask;
  wire       [63:0]   vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_data;
  wire                vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_corrupt;
  reg                 vexiis_0_lsuL1Bus_bus_a_s2mPipe_rValid;
  reg        [2:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode;
  reg        [2:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_param;
  reg        [0:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_source;
  reg        [31:0]   vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_address;
  reg        [2:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_size;
  reg        [7:0]    vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_mask;
  reg        [63:0]   vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_data;
  reg                 vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_corrupt;
  wire                when_Stream_l399_2;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_valid;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_source;
  wire       [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_size;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_denied;
  wire       [63:0]   vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_data;
  wire                vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_corrupt;
  (* keep , syn_keep *) reg                 vexiis_0_lsuL1Bus_noDecoder_toDown_d_rValid /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_param /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [0:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_source /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [2:0]    vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_size /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg                 vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_denied /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [63:0]   vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_data /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg                 vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_corrupt /* synthesis syn_keep = 1 */ ;
  wire                when_Stream_l399_3;
  wire                ioBus_bus_a_valid;
  wire                ioBus_bus_a_ready;
  wire       [2:0]    ioBus_bus_a_payload_opcode;
  wire       [2:0]    ioBus_bus_a_payload_param;
  wire       [31:0]   ioBus_bus_a_payload_address;
  wire       [1:0]    ioBus_bus_a_payload_size;
  wire       [3:0]    ioBus_bus_a_payload_mask;
  wire       [31:0]   ioBus_bus_a_payload_data;
  wire                ioBus_bus_a_payload_corrupt;
  wire                ioBus_bus_d_valid;
  wire                ioBus_bus_d_ready;
  wire       [2:0]    ioBus_bus_d_payload_opcode;
  wire       [2:0]    ioBus_bus_d_payload_param;
  wire       [1:0]    ioBus_bus_d_payload_size;
  wire                ioBus_bus_d_payload_denied;
  wire       [31:0]   ioBus_bus_d_payload_data;
  wire                ioBus_bus_d_payload_corrupt;
  wire                vexiis_0_dBus_to_ioBus_down_bus_a_valid;
  wire                vexiis_0_dBus_to_ioBus_down_bus_a_ready;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_down_bus_a_payload_param;
  wire       [31:0]   vexiis_0_dBus_to_ioBus_down_bus_a_payload_address;
  wire       [1:0]    vexiis_0_dBus_to_ioBus_down_bus_a_payload_size;
  wire       [3:0]    vexiis_0_dBus_to_ioBus_down_bus_a_payload_mask;
  wire       [31:0]   vexiis_0_dBus_to_ioBus_down_bus_a_payload_data;
  wire                vexiis_0_dBus_to_ioBus_down_bus_a_payload_corrupt;
  wire                vexiis_0_dBus_to_ioBus_down_bus_d_valid;
  wire                vexiis_0_dBus_to_ioBus_down_bus_d_ready;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_down_bus_d_payload_param;
  wire       [1:0]    vexiis_0_dBus_to_ioBus_down_bus_d_payload_size;
  wire                vexiis_0_dBus_to_ioBus_down_bus_d_payload_denied;
  wire       [31:0]   vexiis_0_dBus_to_ioBus_down_bus_d_payload_data;
  wire                vexiis_0_dBus_to_ioBus_down_bus_d_payload_corrupt;
  wire                vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_valid;
  wire                vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_ready;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_param;
  wire       [31:0]   vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_address;
  wire       [1:0]    vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_size;
  wire       [3:0]    vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_mask;
  wire       [31:0]   vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_data;
  wire                vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_corrupt;
  reg                 vexiis_0_dBus_to_ioBus_down_bus_a_rValid;
  wire                vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_fire;
  reg        [2:0]    vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode;
  reg        [2:0]    vexiis_0_dBus_to_ioBus_down_bus_a_rData_param;
  reg        [31:0]   vexiis_0_dBus_to_ioBus_down_bus_a_rData_address;
  reg        [1:0]    vexiis_0_dBus_to_ioBus_down_bus_a_rData_size;
  reg        [3:0]    vexiis_0_dBus_to_ioBus_down_bus_a_rData_mask;
  reg        [31:0]   vexiis_0_dBus_to_ioBus_down_bus_a_rData_data;
  reg                 vexiis_0_dBus_to_ioBus_down_bus_a_rData_corrupt;
  wire                ioBus_bus_d_combStage_valid;
  wire                ioBus_bus_d_combStage_ready;
  wire       [2:0]    ioBus_bus_d_combStage_payload_opcode;
  wire       [2:0]    ioBus_bus_d_combStage_payload_param;
  wire       [1:0]    ioBus_bus_d_combStage_payload_size;
  wire                ioBus_bus_d_combStage_payload_denied;
  wire       [31:0]   ioBus_bus_d_combStage_payload_data;
  wire                ioBus_bus_d_combStage_payload_corrupt;
  wire                ioBus_noDecoder_toDown_a_valid;
  wire                ioBus_noDecoder_toDown_a_ready;
  wire       [2:0]    ioBus_noDecoder_toDown_a_payload_opcode;
  wire       [2:0]    ioBus_noDecoder_toDown_a_payload_param;
  wire       [31:0]   ioBus_noDecoder_toDown_a_payload_address;
  wire       [1:0]    ioBus_noDecoder_toDown_a_payload_size;
  wire       [3:0]    ioBus_noDecoder_toDown_a_payload_mask;
  wire       [31:0]   ioBus_noDecoder_toDown_a_payload_data;
  wire                ioBus_noDecoder_toDown_a_payload_corrupt;
  wire                ioBus_noDecoder_toDown_d_valid;
  wire                ioBus_noDecoder_toDown_d_ready;
  wire       [2:0]    ioBus_noDecoder_toDown_d_payload_opcode;
  wire       [2:0]    ioBus_noDecoder_toDown_d_payload_param;
  wire       [1:0]    ioBus_noDecoder_toDown_d_payload_size;
  wire                ioBus_noDecoder_toDown_d_payload_denied;
  wire       [31:0]   ioBus_noDecoder_toDown_d_payload_data;
  wire                ioBus_noDecoder_toDown_d_payload_corrupt;
  wire                splited_mBus_bus_a_valid;
  wire                splited_mBus_bus_a_ready;
  wire       [2:0]    splited_mBus_bus_a_payload_opcode;
  wire       [2:0]    splited_mBus_bus_a_payload_param;
  wire       [1:0]    splited_mBus_bus_a_payload_source;
  wire       [31:0]   splited_mBus_bus_a_payload_address;
  wire       [2:0]    splited_mBus_bus_a_payload_size;
  wire       [7:0]    splited_mBus_bus_a_payload_mask;
  wire       [63:0]   splited_mBus_bus_a_payload_data;
  wire                splited_mBus_bus_a_payload_corrupt;
  wire                splited_mBus_bus_d_valid;
  wire                splited_mBus_bus_d_ready;
  wire       [2:0]    splited_mBus_bus_d_payload_opcode;
  wire       [2:0]    splited_mBus_bus_d_payload_param;
  wire       [1:0]    splited_mBus_bus_d_payload_source;
  wire       [2:0]    splited_mBus_bus_d_payload_size;
  wire                splited_mBus_bus_d_payload_denied;
  wire       [63:0]   splited_mBus_bus_d_payload_data;
  wire                splited_mBus_bus_d_payload_corrupt;
  wire                vexiis_0_iBus_to_splited_mBus_down_bus_a_valid;
  wire                vexiis_0_iBus_to_splited_mBus_down_bus_a_ready;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_param;
  wire       [31:0]   vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_address;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_size;
  wire                vexiis_0_iBus_to_splited_mBus_down_bus_d_valid;
  wire                vexiis_0_iBus_to_splited_mBus_down_bus_d_ready;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_param;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_size;
  wire                vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_denied;
  wire       [63:0]   vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_data;
  wire                vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_corrupt;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_valid;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_source;
  wire       [31:0]   vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_address;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_size;
  wire       [7:0]    vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_mask;
  wire       [63:0]   vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_data;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_corrupt;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_valid;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_source;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_size;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_denied;
  wire       [63:0]   vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_data;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_corrupt;
  wire                peripheral_bus_bus_a_valid;
  wire                peripheral_bus_bus_a_ready;
  wire       [2:0]    peripheral_bus_bus_a_payload_opcode;
  wire       [2:0]    peripheral_bus_bus_a_payload_param;
  wire       [2:0]    peripheral_bus_bus_a_payload_source;
  wire       [31:0]   peripheral_bus_bus_a_payload_address;
  wire       [2:0]    peripheral_bus_bus_a_payload_size;
  wire       [3:0]    peripheral_bus_bus_a_payload_mask;
  wire       [31:0]   peripheral_bus_bus_a_payload_data;
  wire                peripheral_bus_bus_a_payload_corrupt;
  wire                peripheral_bus_bus_d_valid;
  wire                peripheral_bus_bus_d_ready;
  wire       [2:0]    peripheral_bus_bus_d_payload_opcode;
  wire       [2:0]    peripheral_bus_bus_d_payload_param;
  wire       [2:0]    peripheral_bus_bus_d_payload_source;
  wire       [2:0]    peripheral_bus_bus_d_payload_size;
  wire                peripheral_bus_bus_d_payload_denied;
  wire       [31:0]   peripheral_bus_bus_d_payload_data;
  wire                peripheral_bus_bus_d_payload_corrupt;
  wire                ioBus_to_peripheral_bus_down_bus_a_valid;
  wire                ioBus_to_peripheral_bus_down_bus_a_ready;
  wire       [2:0]    ioBus_to_peripheral_bus_down_bus_a_payload_opcode;
  wire       [2:0]    ioBus_to_peripheral_bus_down_bus_a_payload_param;
  wire       [31:0]   ioBus_to_peripheral_bus_down_bus_a_payload_address;
  wire       [1:0]    ioBus_to_peripheral_bus_down_bus_a_payload_size;
  wire       [3:0]    ioBus_to_peripheral_bus_down_bus_a_payload_mask;
  wire       [31:0]   ioBus_to_peripheral_bus_down_bus_a_payload_data;
  wire                ioBus_to_peripheral_bus_down_bus_a_payload_corrupt;
  wire                ioBus_to_peripheral_bus_down_bus_d_valid;
  wire                ioBus_to_peripheral_bus_down_bus_d_ready;
  wire       [2:0]    ioBus_to_peripheral_bus_down_bus_d_payload_opcode;
  wire       [2:0]    ioBus_to_peripheral_bus_down_bus_d_payload_param;
  wire       [1:0]    ioBus_to_peripheral_bus_down_bus_d_payload_size;
  wire                ioBus_to_peripheral_bus_down_bus_d_payload_denied;
  wire       [31:0]   ioBus_to_peripheral_bus_down_bus_d_payload_data;
  wire                ioBus_to_peripheral_bus_down_bus_d_payload_corrupt;
  wire                splited_mBus_to_peripheral_bus_down_bus_a_valid;
  wire                splited_mBus_to_peripheral_bus_down_bus_a_ready;
  wire       [2:0]    splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode;
  wire       [2:0]    splited_mBus_to_peripheral_bus_down_bus_a_payload_param;
  wire       [1:0]    splited_mBus_to_peripheral_bus_down_bus_a_payload_source;
  wire       [31:0]   splited_mBus_to_peripheral_bus_down_bus_a_payload_address;
  wire       [2:0]    splited_mBus_to_peripheral_bus_down_bus_a_payload_size;
  wire       [3:0]    splited_mBus_to_peripheral_bus_down_bus_a_payload_mask;
  wire       [31:0]   splited_mBus_to_peripheral_bus_down_bus_a_payload_data;
  wire                splited_mBus_to_peripheral_bus_down_bus_a_payload_corrupt;
  wire                splited_mBus_to_peripheral_bus_down_bus_d_valid;
  wire                splited_mBus_to_peripheral_bus_down_bus_d_ready;
  wire       [2:0]    splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode;
  wire       [2:0]    splited_mBus_to_peripheral_bus_down_bus_d_payload_param;
  wire       [1:0]    splited_mBus_to_peripheral_bus_down_bus_d_payload_source;
  wire       [2:0]    splited_mBus_to_peripheral_bus_down_bus_d_payload_size;
  wire                splited_mBus_to_peripheral_bus_down_bus_d_payload_denied;
  wire       [31:0]   splited_mBus_to_peripheral_bus_down_bus_d_payload_data;
  wire                splited_mBus_to_peripheral_bus_down_bus_d_payload_corrupt;
  wire                vexiis_0_dBus_to_ioBus_up_bus_a_valid;
  wire                vexiis_0_dBus_to_ioBus_up_bus_a_ready;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_up_bus_a_payload_param;
  wire       [31:0]   vexiis_0_dBus_to_ioBus_up_bus_a_payload_address;
  wire       [1:0]    vexiis_0_dBus_to_ioBus_up_bus_a_payload_size;
  wire       [3:0]    vexiis_0_dBus_to_ioBus_up_bus_a_payload_mask;
  wire       [31:0]   vexiis_0_dBus_to_ioBus_up_bus_a_payload_data;
  wire                vexiis_0_dBus_to_ioBus_up_bus_a_payload_corrupt;
  wire                vexiis_0_dBus_to_ioBus_up_bus_d_valid;
  wire                vexiis_0_dBus_to_ioBus_up_bus_d_ready;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode;
  wire       [2:0]    vexiis_0_dBus_to_ioBus_up_bus_d_payload_param;
  wire       [1:0]    vexiis_0_dBus_to_ioBus_up_bus_d_payload_size;
  wire                vexiis_0_dBus_to_ioBus_up_bus_d_payload_denied;
  wire       [31:0]   vexiis_0_dBus_to_ioBus_up_bus_d_payload_data;
  wire                vexiis_0_dBus_to_ioBus_up_bus_d_payload_corrupt;
  wire                mem_toAxi4_up_bus_a_valid;
  wire                mem_toAxi4_up_bus_a_ready;
  wire       [2:0]    mem_toAxi4_up_bus_a_payload_opcode;
  wire       [2:0]    mem_toAxi4_up_bus_a_payload_param;
  wire       [1:0]    mem_toAxi4_up_bus_a_payload_source;
  wire       [31:0]   mem_toAxi4_up_bus_a_payload_address;
  wire       [2:0]    mem_toAxi4_up_bus_a_payload_size;
  wire       [15:0]   mem_toAxi4_up_bus_a_payload_mask;
  wire       [127:0]  mem_toAxi4_up_bus_a_payload_data;
  wire                mem_toAxi4_up_bus_a_payload_corrupt;
  wire                mem_toAxi4_up_bus_d_valid;
  wire                mem_toAxi4_up_bus_d_ready;
  wire       [2:0]    mem_toAxi4_up_bus_d_payload_opcode;
  wire       [2:0]    mem_toAxi4_up_bus_d_payload_param;
  wire       [1:0]    mem_toAxi4_up_bus_d_payload_source;
  wire       [2:0]    mem_toAxi4_up_bus_d_payload_size;
  wire                mem_toAxi4_up_bus_d_payload_denied;
  wire       [127:0]  mem_toAxi4_up_bus_d_payload_data;
  wire                mem_toAxi4_up_bus_d_payload_corrupt;
  wire                splited_mBus_to_mem_toAxi4_up_down_bus_a_valid;
  wire                splited_mBus_to_mem_toAxi4_up_down_bus_a_ready;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_param;
  wire       [1:0]    splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_source;
  wire       [31:0]   splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_address;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_size;
  wire       [15:0]   splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_mask;
  wire       [127:0]  splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_data;
  wire                splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_corrupt;
  wire                splited_mBus_to_mem_toAxi4_up_down_bus_d_valid;
  wire                splited_mBus_to_mem_toAxi4_up_down_bus_d_ready;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_param;
  wire       [1:0]    splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_source;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_size;
  wire                splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_denied;
  wire       [127:0]  splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_data;
  wire                splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_corrupt;
  wire                vexiis_0_iBus_to_splited_mBus_up_bus_a_valid;
  wire                vexiis_0_iBus_to_splited_mBus_up_bus_a_ready;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_param;
  wire       [31:0]   vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_address;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_size;
  wire                vexiis_0_iBus_to_splited_mBus_up_bus_d_valid;
  wire                vexiis_0_iBus_to_splited_mBus_up_bus_d_ready;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_param;
  wire       [2:0]    vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_size;
  wire                vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_denied;
  wire       [63:0]   vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_data;
  wire                vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_corrupt;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_valid;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_source;
  wire       [31:0]   vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_address;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_size;
  wire       [7:0]    vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_mask;
  wire       [63:0]   vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_data;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_corrupt;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_valid;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_ready;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_param;
  wire       [0:0]    vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_source;
  wire       [2:0]    vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_size;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_denied;
  wire       [63:0]   vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_data;
  wire                vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_corrupt;
  wire                mem_toAxi4_down_aw_valid;
  wire                mem_toAxi4_down_aw_ready;
  wire       [31:0]   mem_toAxi4_down_aw_payload_addr;
  wire       [1:0]    mem_toAxi4_down_aw_payload_id;
  wire       [7:0]    mem_toAxi4_down_aw_payload_len;
  wire       [2:0]    mem_toAxi4_down_aw_payload_size;
  wire       [1:0]    mem_toAxi4_down_aw_payload_burst;
  wire                mem_toAxi4_down_aw_payload_allStrb;
  wire                mem_toAxi4_down_w_valid;
  wire                mem_toAxi4_down_w_ready;
  wire       [127:0]  mem_toAxi4_down_w_payload_data;
  wire       [15:0]   mem_toAxi4_down_w_payload_strb;
  wire                mem_toAxi4_down_w_payload_last;
  wire                mem_toAxi4_down_b_valid;
  wire                mem_toAxi4_down_b_ready;
  wire       [1:0]    mem_toAxi4_down_b_payload_id;
  wire       [1:0]    mem_toAxi4_down_b_payload_resp;
  wire                mem_toAxi4_down_ar_valid;
  wire                mem_toAxi4_down_ar_ready;
  wire       [31:0]   mem_toAxi4_down_ar_payload_addr;
  wire       [1:0]    mem_toAxi4_down_ar_payload_id;
  wire       [7:0]    mem_toAxi4_down_ar_payload_len;
  wire       [2:0]    mem_toAxi4_down_ar_payload_size;
  wire       [1:0]    mem_toAxi4_down_ar_payload_burst;
  wire                mem_toAxi4_down_r_valid;
  wire                mem_toAxi4_down_r_ready;
  wire       [127:0]  mem_toAxi4_down_r_payload_data;
  wire       [1:0]    mem_toAxi4_down_r_payload_id;
  wire       [1:0]    mem_toAxi4_down_r_payload_resp;
  wire                mem_toAxi4_down_r_payload_last;
  wire                peripheral_clint_node_bus_a_valid;
  wire                peripheral_clint_node_bus_a_ready;
  wire       [2:0]    peripheral_clint_node_bus_a_payload_opcode;
  wire       [2:0]    peripheral_clint_node_bus_a_payload_param;
  wire       [2:0]    peripheral_clint_node_bus_a_payload_source;
  wire       [15:0]   peripheral_clint_node_bus_a_payload_address;
  wire       [2:0]    peripheral_clint_node_bus_a_payload_size;
  wire       [3:0]    peripheral_clint_node_bus_a_payload_mask;
  wire       [31:0]   peripheral_clint_node_bus_a_payload_data;
  wire                peripheral_clint_node_bus_a_payload_corrupt;
  wire                peripheral_clint_node_bus_d_valid;
  wire                peripheral_clint_node_bus_d_ready;
  wire       [2:0]    peripheral_clint_node_bus_d_payload_opcode;
  wire       [2:0]    peripheral_clint_node_bus_d_payload_param;
  wire       [2:0]    peripheral_clint_node_bus_d_payload_source;
  wire       [2:0]    peripheral_clint_node_bus_d_payload_size;
  wire                peripheral_clint_node_bus_d_payload_denied;
  wire       [31:0]   peripheral_clint_node_bus_d_payload_data;
  wire                peripheral_clint_node_bus_d_payload_corrupt;
  wire                peripheral_bus_to_peripheral_clint_node_down_bus_a_valid;
  wire                peripheral_bus_to_peripheral_clint_node_down_bus_a_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_source;
  wire       [15:0]   peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_address;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_size;
  wire       [3:0]    peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_mask;
  wire       [31:0]   peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_data;
  wire                peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_corrupt;
  wire                peripheral_bus_to_peripheral_clint_node_down_bus_d_valid;
  wire                peripheral_bus_to_peripheral_clint_node_down_bus_d_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_source;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_size;
  wire                peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_denied;
  wire       [31:0]   peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_data;
  wire                peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_corrupt;
  wire                peripheral_plic_node_bus_a_valid;
  wire                peripheral_plic_node_bus_a_ready;
  wire       [2:0]    peripheral_plic_node_bus_a_payload_opcode;
  wire       [2:0]    peripheral_plic_node_bus_a_payload_param;
  wire       [2:0]    peripheral_plic_node_bus_a_payload_source;
  wire       [21:0]   peripheral_plic_node_bus_a_payload_address;
  wire       [1:0]    peripheral_plic_node_bus_a_payload_size;
  wire       [3:0]    peripheral_plic_node_bus_a_payload_mask;
  wire       [31:0]   peripheral_plic_node_bus_a_payload_data;
  wire                peripheral_plic_node_bus_a_payload_corrupt;
  wire                peripheral_plic_node_bus_d_valid;
  wire                peripheral_plic_node_bus_d_ready;
  wire       [2:0]    peripheral_plic_node_bus_d_payload_opcode;
  wire       [2:0]    peripheral_plic_node_bus_d_payload_param;
  wire       [2:0]    peripheral_plic_node_bus_d_payload_source;
  wire       [1:0]    peripheral_plic_node_bus_d_payload_size;
  wire                peripheral_plic_node_bus_d_payload_denied;
  wire       [31:0]   peripheral_plic_node_bus_d_payload_data;
  wire                peripheral_plic_node_bus_d_payload_corrupt;
  wire                peripheral_bus_to_peripheral_plic_node_down_bus_a_valid;
  wire                peripheral_bus_to_peripheral_plic_node_down_bus_a_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_source;
  wire       [21:0]   peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_address;
  wire       [1:0]    peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_size;
  wire       [3:0]    peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_mask;
  wire       [31:0]   peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_data;
  wire                peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_corrupt;
  wire                peripheral_bus_to_peripheral_plic_node_down_bus_d_valid;
  wire                peripheral_bus_to_peripheral_plic_node_down_bus_d_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_source;
  wire       [1:0]    peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_size;
  wire                peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_denied;
  wire       [31:0]   peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_data;
  wire                peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_corrupt;
  wire                peripheral_toAxiLite4_up_bus_a_valid;
  wire                peripheral_toAxiLite4_up_bus_a_ready;
  wire       [2:0]    peripheral_toAxiLite4_up_bus_a_payload_opcode;
  wire       [2:0]    peripheral_toAxiLite4_up_bus_a_payload_param;
  wire       [2:0]    peripheral_toAxiLite4_up_bus_a_payload_source;
  wire       [31:0]   peripheral_toAxiLite4_up_bus_a_payload_address;
  wire       [2:0]    peripheral_toAxiLite4_up_bus_a_payload_size;
  wire       [3:0]    peripheral_toAxiLite4_up_bus_a_payload_mask;
  wire       [31:0]   peripheral_toAxiLite4_up_bus_a_payload_data;
  wire                peripheral_toAxiLite4_up_bus_a_payload_corrupt;
  wire                peripheral_toAxiLite4_up_bus_d_valid;
  wire                peripheral_toAxiLite4_up_bus_d_ready;
  wire       [2:0]    peripheral_toAxiLite4_up_bus_d_payload_opcode;
  wire       [2:0]    peripheral_toAxiLite4_up_bus_d_payload_param;
  wire       [2:0]    peripheral_toAxiLite4_up_bus_d_payload_source;
  wire       [2:0]    peripheral_toAxiLite4_up_bus_d_payload_size;
  wire                peripheral_toAxiLite4_up_bus_d_payload_denied;
  wire       [31:0]   peripheral_toAxiLite4_up_bus_d_payload_data;
  wire                peripheral_toAxiLite4_up_bus_d_payload_corrupt;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_valid;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_source;
  wire       [31:0]   peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_address;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_size;
  wire       [3:0]    peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_mask;
  wire       [31:0]   peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_data;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_corrupt;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_valid;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_source;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_size;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_denied;
  wire       [31:0]   peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_data;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_corrupt;
  wire                ioBus_to_peripheral_bus_up_bus_a_valid;
  wire                ioBus_to_peripheral_bus_up_bus_a_ready;
  wire       [2:0]    ioBus_to_peripheral_bus_up_bus_a_payload_opcode;
  wire       [2:0]    ioBus_to_peripheral_bus_up_bus_a_payload_param;
  wire       [31:0]   ioBus_to_peripheral_bus_up_bus_a_payload_address;
  wire       [1:0]    ioBus_to_peripheral_bus_up_bus_a_payload_size;
  wire       [3:0]    ioBus_to_peripheral_bus_up_bus_a_payload_mask;
  wire       [31:0]   ioBus_to_peripheral_bus_up_bus_a_payload_data;
  wire                ioBus_to_peripheral_bus_up_bus_a_payload_corrupt;
  wire                ioBus_to_peripheral_bus_up_bus_d_valid;
  wire                ioBus_to_peripheral_bus_up_bus_d_ready;
  wire       [2:0]    ioBus_to_peripheral_bus_up_bus_d_payload_opcode;
  wire       [2:0]    ioBus_to_peripheral_bus_up_bus_d_payload_param;
  wire       [1:0]    ioBus_to_peripheral_bus_up_bus_d_payload_size;
  wire                ioBus_to_peripheral_bus_up_bus_d_payload_denied;
  wire       [31:0]   ioBus_to_peripheral_bus_up_bus_d_payload_data;
  wire                ioBus_to_peripheral_bus_up_bus_d_payload_corrupt;
  wire                splited_mBus_to_mem_toAxi4_up_up_bus_a_valid;
  wire                splited_mBus_to_mem_toAxi4_up_up_bus_a_ready;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_param;
  wire       [1:0]    splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_source;
  wire       [31:0]   splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_address;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_size;
  wire       [7:0]    splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_mask;
  wire       [63:0]   splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_data;
  wire                splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_corrupt;
  wire                splited_mBus_to_mem_toAxi4_up_up_bus_d_valid;
  wire                splited_mBus_to_mem_toAxi4_up_up_bus_d_ready;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_param;
  wire       [1:0]    splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_source;
  wire       [2:0]    splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_size;
  wire                splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_denied;
  wire       [63:0]   splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_data;
  wire                splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_corrupt;
  wire                splited_mBus_to_peripheral_bus_up_bus_a_valid;
  wire                splited_mBus_to_peripheral_bus_up_bus_a_ready;
  wire       [2:0]    splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode;
  wire       [2:0]    splited_mBus_to_peripheral_bus_up_bus_a_payload_param;
  wire       [1:0]    splited_mBus_to_peripheral_bus_up_bus_a_payload_source;
  wire       [31:0]   splited_mBus_to_peripheral_bus_up_bus_a_payload_address;
  wire       [2:0]    splited_mBus_to_peripheral_bus_up_bus_a_payload_size;
  wire       [7:0]    splited_mBus_to_peripheral_bus_up_bus_a_payload_mask;
  wire       [63:0]   splited_mBus_to_peripheral_bus_up_bus_a_payload_data;
  wire                splited_mBus_to_peripheral_bus_up_bus_a_payload_corrupt;
  wire                splited_mBus_to_peripheral_bus_up_bus_d_valid;
  wire                splited_mBus_to_peripheral_bus_up_bus_d_ready;
  wire       [2:0]    splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode;
  wire       [2:0]    splited_mBus_to_peripheral_bus_up_bus_d_payload_param;
  wire       [1:0]    splited_mBus_to_peripheral_bus_up_bus_d_payload_source;
  wire       [2:0]    splited_mBus_to_peripheral_bus_up_bus_d_payload_size;
  wire                splited_mBus_to_peripheral_bus_up_bus_d_payload_denied;
  wire       [63:0]   splited_mBus_to_peripheral_bus_up_bus_d_payload_data;
  wire                splited_mBus_to_peripheral_bus_up_bus_d_payload_corrupt;
  wire                mBusAxi_aw_valid;
  wire                mBusAxi_aw_ready;
  wire       [31:0]   mBusAxi_aw_payload_addr;
  wire       [7:0]    mBusAxi_aw_payload_id;
  wire       [7:0]    mBusAxi_aw_payload_len;
  wire       [2:0]    mBusAxi_aw_payload_size;
  wire       [1:0]    mBusAxi_aw_payload_burst;
  wire                mBusAxi_aw_payload_allStrb;
  wire                mBusAxi_w_valid;
  wire                mBusAxi_w_ready;
  wire       [127:0]  mBusAxi_w_payload_data;
  wire       [15:0]   mBusAxi_w_payload_strb;
  wire                mBusAxi_w_payload_last;
  wire                mBusAxi_b_valid;
  wire                mBusAxi_b_ready;
  wire       [7:0]    mBusAxi_b_payload_id;
  wire       [1:0]    mBusAxi_b_payload_resp;
  wire                mBusAxi_ar_valid;
  wire                mBusAxi_ar_ready;
  wire       [31:0]   mBusAxi_ar_payload_addr;
  wire       [7:0]    mBusAxi_ar_payload_id;
  wire       [7:0]    mBusAxi_ar_payload_len;
  wire       [2:0]    mBusAxi_ar_payload_size;
  wire       [1:0]    mBusAxi_ar_payload_burst;
  wire                mBusAxi_r_valid;
  wire                mBusAxi_r_ready;
  wire       [127:0]  mBusAxi_r_payload_data;
  wire       [7:0]    mBusAxi_r_payload_id;
  wire       [1:0]    mBusAxi_r_payload_resp;
  wire                mBusAxi_r_payload_last;
  wire                mBusAxi_aw_s2mPipe_valid;
  reg                 mBusAxi_aw_s2mPipe_ready;
  wire       [31:0]   mBusAxi_aw_s2mPipe_payload_addr;
  wire       [7:0]    mBusAxi_aw_s2mPipe_payload_id;
  wire       [7:0]    mBusAxi_aw_s2mPipe_payload_len;
  wire       [2:0]    mBusAxi_aw_s2mPipe_payload_size;
  wire       [1:0]    mBusAxi_aw_s2mPipe_payload_burst;
  wire                mBusAxi_aw_s2mPipe_payload_allStrb;
  reg                 mBusAxi_aw_rValidN;
  reg        [31:0]   mBusAxi_aw_rData_addr;
  reg        [7:0]    mBusAxi_aw_rData_id;
  reg        [7:0]    mBusAxi_aw_rData_len;
  reg        [2:0]    mBusAxi_aw_rData_size;
  reg        [1:0]    mBusAxi_aw_rData_burst;
  reg                 mBusAxi_aw_rData_allStrb;
  wire                mBusAxi_aw_s2mPipe_m2sPipe_valid;
  wire                mBusAxi_aw_s2mPipe_m2sPipe_ready;
  wire       [31:0]   mBusAxi_aw_s2mPipe_m2sPipe_payload_addr;
  wire       [7:0]    mBusAxi_aw_s2mPipe_m2sPipe_payload_id;
  wire       [7:0]    mBusAxi_aw_s2mPipe_m2sPipe_payload_len;
  wire       [2:0]    mBusAxi_aw_s2mPipe_m2sPipe_payload_size;
  wire       [1:0]    mBusAxi_aw_s2mPipe_m2sPipe_payload_burst;
  wire                mBusAxi_aw_s2mPipe_m2sPipe_payload_allStrb;
  reg                 mBusAxi_aw_s2mPipe_rValid;
  reg        [31:0]   mBusAxi_aw_s2mPipe_rData_addr;
  reg        [7:0]    mBusAxi_aw_s2mPipe_rData_id;
  reg        [7:0]    mBusAxi_aw_s2mPipe_rData_len;
  reg        [2:0]    mBusAxi_aw_s2mPipe_rData_size;
  reg        [1:0]    mBusAxi_aw_s2mPipe_rData_burst;
  reg                 mBusAxi_aw_s2mPipe_rData_allStrb;
  wire                when_Stream_l399_4;
  wire                mBusAxi_w_s2mPipe_valid;
  reg                 mBusAxi_w_s2mPipe_ready;
  wire       [127:0]  mBusAxi_w_s2mPipe_payload_data;
  wire       [15:0]   mBusAxi_w_s2mPipe_payload_strb;
  wire                mBusAxi_w_s2mPipe_payload_last;
  reg                 mBusAxi_w_rValidN;
  reg        [127:0]  mBusAxi_w_rData_data;
  reg        [15:0]   mBusAxi_w_rData_strb;
  reg                 mBusAxi_w_rData_last;
  wire                mBusAxi_w_s2mPipe_m2sPipe_valid;
  wire                mBusAxi_w_s2mPipe_m2sPipe_ready;
  wire       [127:0]  mBusAxi_w_s2mPipe_m2sPipe_payload_data;
  wire       [15:0]   mBusAxi_w_s2mPipe_m2sPipe_payload_strb;
  wire                mBusAxi_w_s2mPipe_m2sPipe_payload_last;
  reg                 mBusAxi_w_s2mPipe_rValid;
  reg        [127:0]  mBusAxi_w_s2mPipe_rData_data;
  reg        [15:0]   mBusAxi_w_s2mPipe_rData_strb;
  reg                 mBusAxi_w_s2mPipe_rData_last;
  wire                when_Stream_l399_5;
  wire                mBus_b_s2mPipe_valid;
  reg                 mBus_b_s2mPipe_ready;
  wire       [7:0]    mBus_b_s2mPipe_payload_id;
  wire       [1:0]    mBus_b_s2mPipe_payload_resp;
  reg                 mBus_b_rValidN;
  reg        [7:0]    mBus_b_rData_id;
  reg        [1:0]    mBus_b_rData_resp;
  wire                mBus_b_s2mPipe_m2sPipe_valid;
  wire                mBus_b_s2mPipe_m2sPipe_ready;
  wire       [7:0]    mBus_b_s2mPipe_m2sPipe_payload_id;
  wire       [1:0]    mBus_b_s2mPipe_m2sPipe_payload_resp;
  reg                 mBus_b_s2mPipe_rValid;
  reg        [7:0]    mBus_b_s2mPipe_rData_id;
  reg        [1:0]    mBus_b_s2mPipe_rData_resp;
  wire                when_Stream_l399_6;
  wire                mBusAxi_ar_s2mPipe_valid;
  reg                 mBusAxi_ar_s2mPipe_ready;
  wire       [31:0]   mBusAxi_ar_s2mPipe_payload_addr;
  wire       [7:0]    mBusAxi_ar_s2mPipe_payload_id;
  wire       [7:0]    mBusAxi_ar_s2mPipe_payload_len;
  wire       [2:0]    mBusAxi_ar_s2mPipe_payload_size;
  wire       [1:0]    mBusAxi_ar_s2mPipe_payload_burst;
  reg                 mBusAxi_ar_rValidN;
  reg        [31:0]   mBusAxi_ar_rData_addr;
  reg        [7:0]    mBusAxi_ar_rData_id;
  reg        [7:0]    mBusAxi_ar_rData_len;
  reg        [2:0]    mBusAxi_ar_rData_size;
  reg        [1:0]    mBusAxi_ar_rData_burst;
  wire                mBusAxi_ar_s2mPipe_m2sPipe_valid;
  wire                mBusAxi_ar_s2mPipe_m2sPipe_ready;
  wire       [31:0]   mBusAxi_ar_s2mPipe_m2sPipe_payload_addr;
  wire       [7:0]    mBusAxi_ar_s2mPipe_m2sPipe_payload_id;
  wire       [7:0]    mBusAxi_ar_s2mPipe_m2sPipe_payload_len;
  wire       [2:0]    mBusAxi_ar_s2mPipe_m2sPipe_payload_size;
  wire       [1:0]    mBusAxi_ar_s2mPipe_m2sPipe_payload_burst;
  reg                 mBusAxi_ar_s2mPipe_rValid;
  reg        [31:0]   mBusAxi_ar_s2mPipe_rData_addr;
  reg        [7:0]    mBusAxi_ar_s2mPipe_rData_id;
  reg        [7:0]    mBusAxi_ar_s2mPipe_rData_len;
  reg        [2:0]    mBusAxi_ar_s2mPipe_rData_size;
  reg        [1:0]    mBusAxi_ar_s2mPipe_rData_burst;
  wire                when_Stream_l399_7;
  wire                mBus_r_s2mPipe_valid;
  reg                 mBus_r_s2mPipe_ready;
  wire       [127:0]  mBus_r_s2mPipe_payload_data;
  wire       [7:0]    mBus_r_s2mPipe_payload_id;
  wire       [1:0]    mBus_r_s2mPipe_payload_resp;
  wire                mBus_r_s2mPipe_payload_last;
  reg                 mBus_r_rValidN;
  reg        [127:0]  mBus_r_rData_data;
  reg        [7:0]    mBus_r_rData_id;
  reg        [1:0]    mBus_r_rData_resp;
  reg                 mBus_r_rData_last;
  wire                mBus_r_s2mPipe_m2sPipe_valid;
  wire                mBus_r_s2mPipe_m2sPipe_ready;
  wire       [127:0]  mBus_r_s2mPipe_m2sPipe_payload_data;
  wire       [7:0]    mBus_r_s2mPipe_m2sPipe_payload_id;
  wire       [1:0]    mBus_r_s2mPipe_m2sPipe_payload_resp;
  wire                mBus_r_s2mPipe_m2sPipe_payload_last;
  reg                 mBus_r_s2mPipe_rValid;
  reg        [127:0]  mBus_r_s2mPipe_rData_data;
  reg        [7:0]    mBus_r_s2mPipe_rData_id;
  reg        [1:0]    mBus_r_s2mPipe_rData_resp;
  reg                 mBus_r_s2mPipe_rData_last;
  wire                when_Stream_l399_8;
  wire                peripheral_toAxiLite4_down_aw_valid;
  wire                peripheral_toAxiLite4_down_aw_ready;
  wire       [31:0]   peripheral_toAxiLite4_down_aw_payload_addr;
  wire       [2:0]    peripheral_toAxiLite4_down_aw_payload_prot;
  wire                peripheral_toAxiLite4_down_w_valid;
  wire                peripheral_toAxiLite4_down_w_ready;
  wire       [31:0]   peripheral_toAxiLite4_down_w_payload_data;
  wire       [3:0]    peripheral_toAxiLite4_down_w_payload_strb;
  wire                peripheral_toAxiLite4_down_b_valid;
  wire                peripheral_toAxiLite4_down_b_ready;
  wire       [1:0]    peripheral_toAxiLite4_down_b_payload_resp;
  wire                peripheral_toAxiLite4_down_ar_valid;
  wire                peripheral_toAxiLite4_down_ar_ready;
  wire       [31:0]   peripheral_toAxiLite4_down_ar_payload_addr;
  wire       [2:0]    peripheral_toAxiLite4_down_ar_payload_prot;
  wire                peripheral_toAxiLite4_down_r_valid;
  wire                peripheral_toAxiLite4_down_r_ready;
  wire       [31:0]   peripheral_toAxiLite4_down_r_payload_data;
  wire       [1:0]    peripheral_toAxiLite4_down_r_payload_resp;
  wire                peripheral_bus_to_peripheral_clint_node_up_bus_a_valid;
  wire                peripheral_bus_to_peripheral_clint_node_up_bus_a_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_source;
  wire       [15:0]   peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_address;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_size;
  wire       [3:0]    peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_mask;
  wire       [31:0]   peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_data;
  wire                peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_corrupt;
  wire                peripheral_bus_to_peripheral_clint_node_up_bus_d_valid;
  wire                peripheral_bus_to_peripheral_clint_node_up_bus_d_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_source;
  wire       [2:0]    peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_size;
  wire                peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_denied;
  wire       [31:0]   peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_data;
  wire                peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_corrupt;
  wire                peripheral_bus_to_peripheral_plic_node_up_bus_a_valid;
  wire                peripheral_bus_to_peripheral_plic_node_up_bus_a_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_source;
  wire       [21:0]   peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_address;
  wire       [1:0]    peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_size;
  wire       [3:0]    peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_mask;
  wire       [31:0]   peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_data;
  wire                peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_corrupt;
  wire                peripheral_bus_to_peripheral_plic_node_up_bus_d_valid;
  wire                peripheral_bus_to_peripheral_plic_node_up_bus_d_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_source;
  wire       [1:0]    peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_size;
  wire                peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_denied;
  wire       [31:0]   peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_data;
  wire                peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_corrupt;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_valid;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_source;
  wire       [31:0]   peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_address;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_size;
  wire       [3:0]    peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_mask;
  wire       [31:0]   peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_data;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_corrupt;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_valid;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_ready;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_param;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_source;
  wire       [2:0]    peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_size;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_denied;
  wire       [31:0]   peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_data;
  wire                peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_corrupt;
  wire                peripheral_bus_bus_a_halfPipe_valid;
  wire                peripheral_bus_bus_a_halfPipe_ready;
  wire       [2:0]    peripheral_bus_bus_a_halfPipe_payload_opcode;
  wire       [2:0]    peripheral_bus_bus_a_halfPipe_payload_param;
  wire       [2:0]    peripheral_bus_bus_a_halfPipe_payload_source;
  wire       [31:0]   peripheral_bus_bus_a_halfPipe_payload_address;
  wire       [2:0]    peripheral_bus_bus_a_halfPipe_payload_size;
  wire       [3:0]    peripheral_bus_bus_a_halfPipe_payload_mask;
  wire       [31:0]   peripheral_bus_bus_a_halfPipe_payload_data;
  wire                peripheral_bus_bus_a_halfPipe_payload_corrupt;
  reg                 peripheral_bus_bus_a_rValid;
  wire                peripheral_bus_bus_a_halfPipe_fire;
  reg        [2:0]    peripheral_bus_bus_a_rData_opcode;
  reg        [2:0]    peripheral_bus_bus_a_rData_param;
  reg        [2:0]    peripheral_bus_bus_a_rData_source;
  reg        [31:0]   peripheral_bus_bus_a_rData_address;
  reg        [2:0]    peripheral_bus_bus_a_rData_size;
  reg        [3:0]    peripheral_bus_bus_a_rData_mask;
  reg        [31:0]   peripheral_bus_bus_a_rData_data;
  reg                 peripheral_bus_bus_a_rData_corrupt;
  wire                io_up_d_halfPipe_valid;
  wire                io_up_d_halfPipe_ready;
  wire       [2:0]    io_up_d_halfPipe_payload_opcode;
  wire       [2:0]    io_up_d_halfPipe_payload_param;
  wire       [2:0]    io_up_d_halfPipe_payload_source;
  wire       [2:0]    io_up_d_halfPipe_payload_size;
  wire                io_up_d_halfPipe_payload_denied;
  wire       [31:0]   io_up_d_halfPipe_payload_data;
  wire                io_up_d_halfPipe_payload_corrupt;
  reg                 io_up_d_rValid;
  wire                io_up_d_halfPipe_fire;
  reg        [2:0]    io_up_d_rData_opcode;
  reg        [2:0]    io_up_d_rData_param;
  reg        [2:0]    io_up_d_rData_source;
  reg        [2:0]    io_up_d_rData_size;
  reg                 io_up_d_rData_denied;
  reg        [31:0]   io_up_d_rData_data;
  reg                 io_up_d_rData_corrupt;
  wire                peripheral_toAxiLite4_down_aw_halfPipe_valid;
  wire                peripheral_toAxiLite4_down_aw_halfPipe_ready;
  wire       [31:0]   peripheral_toAxiLite4_down_aw_halfPipe_payload_addr;
  wire       [2:0]    peripheral_toAxiLite4_down_aw_halfPipe_payload_prot;
  reg                 peripheral_toAxiLite4_down_aw_rValid;
  wire                peripheral_toAxiLite4_down_aw_halfPipe_fire;
  reg        [31:0]   peripheral_toAxiLite4_down_aw_rData_addr;
  reg        [2:0]    peripheral_toAxiLite4_down_aw_rData_prot;
  wire                peripheral_toAxiLite4_down_w_halfPipe_valid;
  wire                peripheral_toAxiLite4_down_w_halfPipe_ready;
  wire       [31:0]   peripheral_toAxiLite4_down_w_halfPipe_payload_data;
  wire       [3:0]    peripheral_toAxiLite4_down_w_halfPipe_payload_strb;
  reg                 peripheral_toAxiLite4_down_w_rValid;
  wire                peripheral_toAxiLite4_down_w_halfPipe_fire;
  reg        [31:0]   peripheral_toAxiLite4_down_w_rData_data;
  reg        [3:0]    peripheral_toAxiLite4_down_w_rData_strb;
  wire                pBus_b_halfPipe_valid;
  wire                pBus_b_halfPipe_ready;
  wire       [1:0]    pBus_b_halfPipe_payload_resp;
  reg                 pBus_b_rValid;
  wire                pBus_b_halfPipe_fire;
  reg        [1:0]    pBus_b_rData_resp;
  wire                peripheral_toAxiLite4_down_ar_halfPipe_valid;
  wire                peripheral_toAxiLite4_down_ar_halfPipe_ready;
  wire       [31:0]   peripheral_toAxiLite4_down_ar_halfPipe_payload_addr;
  wire       [2:0]    peripheral_toAxiLite4_down_ar_halfPipe_payload_prot;
  reg                 peripheral_toAxiLite4_down_ar_rValid;
  wire                peripheral_toAxiLite4_down_ar_halfPipe_fire;
  reg        [31:0]   peripheral_toAxiLite4_down_ar_rData_addr;
  reg        [2:0]    peripheral_toAxiLite4_down_ar_rData_prot;
  wire                pBus_r_halfPipe_valid;
  wire                pBus_r_halfPipe_ready;
  wire       [31:0]   pBus_r_halfPipe_payload_data;
  wire       [1:0]    pBus_r_halfPipe_payload_resp;
  reg                 pBus_r_rValid;
  wire                pBus_r_halfPipe_fire;
  reg        [31:0]   pBus_r_rData_data;
  reg        [1:0]    pBus_r_rData_resp;
  wire       [7:0]    debugIn;
  reg        [7:0]    debugIn_delay_1;
  `ifndef SYNTHESIS
  reg [127:0] vexiis_0_dBus_bus_a_payload_opcode_string;
  reg [119:0] vexiis_0_dBus_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_dBus_noDecoder_toDown_a_payload_opcode_string;
  reg [119:0] vexiis_0_dBus_noDecoder_toDown_d_payload_opcode_string;
  reg [127:0] vexiis_0_dBus_bus_a_halfPipe_payload_opcode_string;
  reg [127:0] vexiis_0_dBus_bus_a_rData_opcode_string;
  reg [119:0] vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode_string;
  reg [119:0] vexiis_0_dBus_noDecoder_toDown_d_rData_opcode_string;
  reg [127:0] vexiis_0_iBus_bus_a_payload_opcode_string;
  reg [119:0] vexiis_0_iBus_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_iBus_noDecoder_toDown_a_payload_opcode_string;
  reg [119:0] vexiis_0_iBus_noDecoder_toDown_d_payload_opcode_string;
  reg [127:0] vexiis_0_iBus_bus_a_halfPipe_payload_opcode_string;
  reg [127:0] vexiis_0_iBus_bus_a_rData_opcode_string;
  reg [127:0] vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode_string;
  reg [127:0] vexiis_0_iBus_bus_a_halfPipe_rData_opcode_string;
  reg [119:0] vexiis_0_iBus_noDecoder_connection_payload_opcode_string;
  reg [119:0] vexiis_0_iBus_noDecoder_toDown_d_rData_opcode_string;
  reg [127:0] vexiis_0_lsuL1Bus_bus_a_payload_opcode_string;
  reg [119:0] vexiis_0_lsuL1Bus_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode_string;
  reg [119:0] vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode_string;
  reg [127:0] vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string;
  reg [127:0] vexiis_0_lsuL1Bus_bus_a_rData_opcode_string;
  reg [127:0] _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string;
  reg [127:0] vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode_string;
  reg [127:0] vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode_string;
  reg [119:0] vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode_string;
  reg [119:0] vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode_string;
  reg [127:0] ioBus_bus_a_payload_opcode_string;
  reg [119:0] ioBus_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode_string;
  reg [119:0] vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode_string;
  reg [127:0] vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode_string;
  reg [119:0] ioBus_bus_d_combStage_payload_opcode_string;
  reg [127:0] ioBus_noDecoder_toDown_a_payload_opcode_string;
  reg [119:0] ioBus_noDecoder_toDown_d_payload_opcode_string;
  reg [127:0] splited_mBus_bus_a_payload_opcode_string;
  reg [119:0] splited_mBus_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode_string;
  reg [119:0] vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode_string;
  reg [119:0] vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode_string;
  reg [127:0] peripheral_bus_bus_a_payload_opcode_string;
  reg [119:0] peripheral_bus_bus_d_payload_opcode_string;
  reg [127:0] ioBus_to_peripheral_bus_down_bus_a_payload_opcode_string;
  reg [119:0] ioBus_to_peripheral_bus_down_bus_d_payload_opcode_string;
  reg [127:0] splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode_string;
  reg [119:0] splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode_string;
  reg [119:0] vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode_string;
  reg [127:0] mem_toAxi4_up_bus_a_payload_opcode_string;
  reg [119:0] mem_toAxi4_up_bus_d_payload_opcode_string;
  reg [127:0] splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode_string;
  reg [119:0] splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode_string;
  reg [119:0] vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode_string;
  reg [127:0] vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode_string;
  reg [119:0] vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode_string;
  reg [127:0] peripheral_clint_node_bus_a_payload_opcode_string;
  reg [119:0] peripheral_clint_node_bus_d_payload_opcode_string;
  reg [127:0] peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode_string;
  reg [119:0] peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode_string;
  reg [127:0] peripheral_plic_node_bus_a_payload_opcode_string;
  reg [119:0] peripheral_plic_node_bus_d_payload_opcode_string;
  reg [127:0] peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode_string;
  reg [119:0] peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode_string;
  reg [127:0] peripheral_toAxiLite4_up_bus_a_payload_opcode_string;
  reg [119:0] peripheral_toAxiLite4_up_bus_d_payload_opcode_string;
  reg [127:0] peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode_string;
  reg [119:0] peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode_string;
  reg [127:0] ioBus_to_peripheral_bus_up_bus_a_payload_opcode_string;
  reg [119:0] ioBus_to_peripheral_bus_up_bus_d_payload_opcode_string;
  reg [127:0] splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode_string;
  reg [119:0] splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode_string;
  reg [127:0] splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode_string;
  reg [119:0] splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode_string;
  reg [127:0] peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode_string;
  reg [119:0] peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode_string;
  reg [127:0] peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode_string;
  reg [119:0] peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode_string;
  reg [127:0] peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode_string;
  reg [119:0] peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode_string;
  reg [127:0] peripheral_bus_bus_a_halfPipe_payload_opcode_string;
  reg [127:0] peripheral_bus_bus_a_rData_opcode_string;
  reg [119:0] io_up_d_halfPipe_payload_opcode_string;
  reg [119:0] io_up_d_rData_opcode_string;
  `endif


  VexiiRiscv vexiis_0_logic_core (
    .CfuPlugin_logic_bus_cmd_valid                         (vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_valid                              ), //o
    .CfuPlugin_logic_bus_cmd_ready                         (vexiis_0_cfuBus_node_cmd_ready                                                 ), //i
    .CfuPlugin_logic_bus_cmd_payload_function_id           (vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_function_id[2:0]           ), //o
    .CfuPlugin_logic_bus_cmd_payload_inputs_0              (vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_inputs_0[31:0]             ), //o
    .CfuPlugin_logic_bus_cmd_payload_inputs_1              (vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_inputs_1[31:0]             ), //o
    .CfuPlugin_logic_bus_cmd_payload_state_index           (vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_state_index[2:0]           ), //o
    .CfuPlugin_logic_bus_cmd_payload_cfu_index             (vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_cfu_index[3:0]             ), //o
    .CfuPlugin_logic_bus_cmd_payload_raw_insn              (vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_raw_insn[31:0]             ), //o
    .CfuPlugin_logic_bus_rsp_valid                         (vexiis_0_cfuBus_node_rsp_valid                                                 ), //i
    .CfuPlugin_logic_bus_rsp_ready                         (vexiis_0_logic_core_CfuPlugin_logic_bus_rsp_ready                              ), //o
    .CfuPlugin_logic_bus_rsp_payload_outputs_0             (vexiis_0_cfuBus_node_rsp_payload_outputs_0[31:0]                               ), //i
    .PrivilegedPlugin_logic_rdtime                         (vexiis_0_priv_rdtime[63:0]                                                     ), //i
    .PrivilegedPlugin_logic_harts_0_int_m_timer            (vexiis_0_priv_mti_flag                                                         ), //i
    .PrivilegedPlugin_logic_harts_0_int_m_software         (vexiis_0_priv_msi_flag                                                         ), //i
    .PrivilegedPlugin_logic_harts_0_int_m_external         (vexiis_0_priv_mei_flag                                                         ), //i
    .PrivilegedPlugin_logic_harts_0_int_s_external         (vexiis_0_priv_sei_flag                                                         ), //i
    .FetchL1TileLinkPlugin_logic_down_a_valid              (vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_valid                   ), //o
    .FetchL1TileLinkPlugin_logic_down_a_ready              (vexiis_0_iBus_bus_a_ready                                                      ), //i
    .FetchL1TileLinkPlugin_logic_down_a_payload_opcode     (vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_opcode[2:0]     ), //o
    .FetchL1TileLinkPlugin_logic_down_a_payload_param      (vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_param[2:0]      ), //o
    .FetchL1TileLinkPlugin_logic_down_a_payload_address    (vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_address[31:0]   ), //o
    .FetchL1TileLinkPlugin_logic_down_a_payload_size       (vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_size[2:0]       ), //o
    .FetchL1TileLinkPlugin_logic_down_d_valid              (vexiis_0_iBus_bus_d_valid                                                      ), //i
    .FetchL1TileLinkPlugin_logic_down_d_ready              (vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_d_ready                   ), //o
    .FetchL1TileLinkPlugin_logic_down_d_payload_opcode     (vexiis_0_iBus_bus_d_payload_opcode[2:0]                                        ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_param      (vexiis_0_iBus_bus_d_payload_param[2:0]                                         ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_size       (vexiis_0_iBus_bus_d_payload_size[2:0]                                          ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_denied     (vexiis_0_iBus_bus_d_payload_denied                                             ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_data       (vexiis_0_iBus_bus_d_payload_data[63:0]                                         ), //i
    .FetchL1TileLinkPlugin_logic_down_d_payload_corrupt    (vexiis_0_iBus_bus_d_payload_corrupt                                            ), //i
    .LsuL1TileLinkPlugin_logic_down_a_valid                (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_valid                     ), //o
    .LsuL1TileLinkPlugin_logic_down_a_ready                (vexiis_0_lsuL1Bus_bus_a_ready                                                  ), //i
    .LsuL1TileLinkPlugin_logic_down_a_payload_opcode       (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_opcode[2:0]       ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_param        (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_param[2:0]        ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_source       (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_source            ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_address      (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_address[31:0]     ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_size         (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_size[2:0]         ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_mask         (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_mask[7:0]         ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_data         (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_data[63:0]        ), //o
    .LsuL1TileLinkPlugin_logic_down_a_payload_corrupt      (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_corrupt           ), //o
    .LsuL1TileLinkPlugin_logic_down_d_valid                (vexiis_0_lsuL1Bus_bus_d_valid                                                  ), //i
    .LsuL1TileLinkPlugin_logic_down_d_ready                (vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_d_ready                     ), //o
    .LsuL1TileLinkPlugin_logic_down_d_payload_opcode       (vexiis_0_lsuL1Bus_bus_d_payload_opcode[2:0]                                    ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_param        (vexiis_0_lsuL1Bus_bus_d_payload_param[2:0]                                     ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_source       (vexiis_0_lsuL1Bus_bus_d_payload_source                                         ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_size         (vexiis_0_lsuL1Bus_bus_d_payload_size[2:0]                                      ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_denied       (vexiis_0_lsuL1Bus_bus_d_payload_denied                                         ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_data         (vexiis_0_lsuL1Bus_bus_d_payload_data[63:0]                                     ), //i
    .LsuL1TileLinkPlugin_logic_down_d_payload_corrupt      (vexiis_0_lsuL1Bus_bus_d_payload_corrupt                                        ), //i
    .LsuTileLinkPlugin_logic_bridge_down_a_valid           (vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_valid                ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_ready           (vexiis_0_dBus_bus_a_ready                                                      ), //i
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode  (vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode[2:0]  ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_param   (vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_param[2:0]   ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_address (vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_address[31:0]), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_size    (vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_size[1:0]    ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_mask    (vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_mask[3:0]    ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_data    (vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_data[31:0]   ), //o
    .LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt (vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt      ), //o
    .LsuTileLinkPlugin_logic_bridge_down_d_valid           (vexiis_0_dBus_bus_d_valid                                                      ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_ready           (vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_d_ready                ), //o
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode  (vexiis_0_dBus_bus_d_payload_opcode[2:0]                                        ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_param   (vexiis_0_dBus_bus_d_payload_param[2:0]                                         ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_size    (vexiis_0_dBus_bus_d_payload_size[1:0]                                          ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_denied  (vexiis_0_dBus_bus_d_payload_denied                                             ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_data    (vexiis_0_dBus_bus_d_payload_data[31:0]                                         ), //i
    .LsuTileLinkPlugin_logic_bridge_down_d_payload_corrupt (vexiis_0_dBus_bus_d_payload_corrupt                                            ), //i
    .litex_clk                                             (litex_clk                                                                      ), //i
    .cpuResetCtrl_reset                                    (cpuResetCtrl_reset                                                             )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC cpuResetCtrl_fiber_aggregator_asyncBuffers_0 (
    .io_dataIn   (1'b0                                                   ), //i
    .io_dataOut  (cpuResetCtrl_fiber_aggregator_asyncBuffers_0_io_dataOut), //o
    .litex_clk   (litex_clk                                              ), //i
    .litex_reset (litex_reset                                            )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_1 cpuResetCtrl_fiber_buffer (
    .io_dataIn                       (1'b0                                ), //i
    .io_dataOut                      (cpuResetCtrl_fiber_buffer_io_dataOut), //o
    .litex_clk                       (litex_clk                           ), //i
    .cpuResetCtrl_fiber_holder_reset (cpuResetCtrl_fiber_holder_reset     )  //i
  );
  Arbiter splited_mBus_arbiter_core (
    .io_ups_0_a_valid           (vexiis_0_iBus_to_splited_mBus_down_bus_a_valid                    ), //i
    .io_ups_0_a_ready           (splited_mBus_arbiter_core_io_ups_0_a_ready                        ), //o
    .io_ups_0_a_payload_opcode  (vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode[2:0]      ), //i
    .io_ups_0_a_payload_param   (vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_param[2:0]       ), //i
    .io_ups_0_a_payload_address (vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_address[31:0]    ), //i
    .io_ups_0_a_payload_size    (vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_size[2:0]        ), //i
    .io_ups_0_d_valid           (splited_mBus_arbiter_core_io_ups_0_d_valid                        ), //o
    .io_ups_0_d_ready           (vexiis_0_iBus_to_splited_mBus_down_bus_d_ready                    ), //i
    .io_ups_0_d_payload_opcode  (splited_mBus_arbiter_core_io_ups_0_d_payload_opcode[2:0]          ), //o
    .io_ups_0_d_payload_param   (splited_mBus_arbiter_core_io_ups_0_d_payload_param[2:0]           ), //o
    .io_ups_0_d_payload_size    (splited_mBus_arbiter_core_io_ups_0_d_payload_size[2:0]            ), //o
    .io_ups_0_d_payload_denied  (splited_mBus_arbiter_core_io_ups_0_d_payload_denied               ), //o
    .io_ups_0_d_payload_data    (splited_mBus_arbiter_core_io_ups_0_d_payload_data[63:0]           ), //o
    .io_ups_0_d_payload_corrupt (splited_mBus_arbiter_core_io_ups_0_d_payload_corrupt              ), //o
    .io_ups_1_a_valid           (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_valid                ), //i
    .io_ups_1_a_ready           (splited_mBus_arbiter_core_io_ups_1_a_ready                        ), //o
    .io_ups_1_a_payload_opcode  (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode[2:0]  ), //i
    .io_ups_1_a_payload_param   (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_param[2:0]   ), //i
    .io_ups_1_a_payload_source  (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_source       ), //i
    .io_ups_1_a_payload_address (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_address[31:0]), //i
    .io_ups_1_a_payload_size    (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_size[2:0]    ), //i
    .io_ups_1_a_payload_mask    (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_mask[7:0]    ), //i
    .io_ups_1_a_payload_data    (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_data[63:0]   ), //i
    .io_ups_1_a_payload_corrupt (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_corrupt      ), //i
    .io_ups_1_d_valid           (splited_mBus_arbiter_core_io_ups_1_d_valid                        ), //o
    .io_ups_1_d_ready           (vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_ready                ), //i
    .io_ups_1_d_payload_opcode  (splited_mBus_arbiter_core_io_ups_1_d_payload_opcode[2:0]          ), //o
    .io_ups_1_d_payload_param   (splited_mBus_arbiter_core_io_ups_1_d_payload_param[2:0]           ), //o
    .io_ups_1_d_payload_source  (splited_mBus_arbiter_core_io_ups_1_d_payload_source               ), //o
    .io_ups_1_d_payload_size    (splited_mBus_arbiter_core_io_ups_1_d_payload_size[2:0]            ), //o
    .io_ups_1_d_payload_denied  (splited_mBus_arbiter_core_io_ups_1_d_payload_denied               ), //o
    .io_ups_1_d_payload_data    (splited_mBus_arbiter_core_io_ups_1_d_payload_data[63:0]           ), //o
    .io_ups_1_d_payload_corrupt (splited_mBus_arbiter_core_io_ups_1_d_payload_corrupt              ), //o
    .io_down_a_valid            (splited_mBus_arbiter_core_io_down_a_valid                         ), //o
    .io_down_a_ready            (splited_mBus_bus_a_ready                                          ), //i
    .io_down_a_payload_opcode   (splited_mBus_arbiter_core_io_down_a_payload_opcode[2:0]           ), //o
    .io_down_a_payload_param    (splited_mBus_arbiter_core_io_down_a_payload_param[2:0]            ), //o
    .io_down_a_payload_source   (splited_mBus_arbiter_core_io_down_a_payload_source[1:0]           ), //o
    .io_down_a_payload_address  (splited_mBus_arbiter_core_io_down_a_payload_address[31:0]         ), //o
    .io_down_a_payload_size     (splited_mBus_arbiter_core_io_down_a_payload_size[2:0]             ), //o
    .io_down_a_payload_mask     (splited_mBus_arbiter_core_io_down_a_payload_mask[7:0]             ), //o
    .io_down_a_payload_data     (splited_mBus_arbiter_core_io_down_a_payload_data[63:0]            ), //o
    .io_down_a_payload_corrupt  (splited_mBus_arbiter_core_io_down_a_payload_corrupt               ), //o
    .io_down_d_valid            (splited_mBus_bus_d_valid                                          ), //i
    .io_down_d_ready            (splited_mBus_arbiter_core_io_down_d_ready                         ), //o
    .io_down_d_payload_opcode   (splited_mBus_bus_d_payload_opcode[2:0]                            ), //i
    .io_down_d_payload_param    (splited_mBus_bus_d_payload_param[2:0]                             ), //i
    .io_down_d_payload_source   (splited_mBus_bus_d_payload_source[1:0]                            ), //i
    .io_down_d_payload_size     (splited_mBus_bus_d_payload_size[2:0]                              ), //i
    .io_down_d_payload_denied   (splited_mBus_bus_d_payload_denied                                 ), //i
    .io_down_d_payload_data     (splited_mBus_bus_d_payload_data[63:0]                             ), //i
    .io_down_d_payload_corrupt  (splited_mBus_bus_d_payload_corrupt                                ), //i
    .litex_clk                  (litex_clk                                                         ), //i
    .cpuResetCtrl_reset         (cpuResetCtrl_reset                                                )  //i
  );
  Arbiter_1 peripheral_bus_arbiter_core (
    .io_ups_0_a_valid           (ioBus_to_peripheral_bus_down_bus_a_valid                       ), //i
    .io_ups_0_a_ready           (peripheral_bus_arbiter_core_io_ups_0_a_ready                   ), //o
    .io_ups_0_a_payload_opcode  (ioBus_to_peripheral_bus_down_bus_a_payload_opcode[2:0]         ), //i
    .io_ups_0_a_payload_param   (ioBus_to_peripheral_bus_down_bus_a_payload_param[2:0]          ), //i
    .io_ups_0_a_payload_address (ioBus_to_peripheral_bus_down_bus_a_payload_address[31:0]       ), //i
    .io_ups_0_a_payload_size    (ioBus_to_peripheral_bus_down_bus_a_payload_size[1:0]           ), //i
    .io_ups_0_a_payload_mask    (ioBus_to_peripheral_bus_down_bus_a_payload_mask[3:0]           ), //i
    .io_ups_0_a_payload_data    (ioBus_to_peripheral_bus_down_bus_a_payload_data[31:0]          ), //i
    .io_ups_0_a_payload_corrupt (ioBus_to_peripheral_bus_down_bus_a_payload_corrupt             ), //i
    .io_ups_0_d_valid           (peripheral_bus_arbiter_core_io_ups_0_d_valid                   ), //o
    .io_ups_0_d_ready           (ioBus_to_peripheral_bus_down_bus_d_ready                       ), //i
    .io_ups_0_d_payload_opcode  (peripheral_bus_arbiter_core_io_ups_0_d_payload_opcode[2:0]     ), //o
    .io_ups_0_d_payload_param   (peripheral_bus_arbiter_core_io_ups_0_d_payload_param[2:0]      ), //o
    .io_ups_0_d_payload_size    (peripheral_bus_arbiter_core_io_ups_0_d_payload_size[1:0]       ), //o
    .io_ups_0_d_payload_denied  (peripheral_bus_arbiter_core_io_ups_0_d_payload_denied          ), //o
    .io_ups_0_d_payload_data    (peripheral_bus_arbiter_core_io_ups_0_d_payload_data[31:0]      ), //o
    .io_ups_0_d_payload_corrupt (peripheral_bus_arbiter_core_io_ups_0_d_payload_corrupt         ), //o
    .io_ups_1_a_valid           (splited_mBus_to_peripheral_bus_down_bus_a_valid                ), //i
    .io_ups_1_a_ready           (peripheral_bus_arbiter_core_io_ups_1_a_ready                   ), //o
    .io_ups_1_a_payload_opcode  (splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode[2:0]  ), //i
    .io_ups_1_a_payload_param   (splited_mBus_to_peripheral_bus_down_bus_a_payload_param[2:0]   ), //i
    .io_ups_1_a_payload_source  (splited_mBus_to_peripheral_bus_down_bus_a_payload_source[1:0]  ), //i
    .io_ups_1_a_payload_address (splited_mBus_to_peripheral_bus_down_bus_a_payload_address[31:0]), //i
    .io_ups_1_a_payload_size    (splited_mBus_to_peripheral_bus_down_bus_a_payload_size[2:0]    ), //i
    .io_ups_1_a_payload_mask    (splited_mBus_to_peripheral_bus_down_bus_a_payload_mask[3:0]    ), //i
    .io_ups_1_a_payload_data    (splited_mBus_to_peripheral_bus_down_bus_a_payload_data[31:0]   ), //i
    .io_ups_1_a_payload_corrupt (splited_mBus_to_peripheral_bus_down_bus_a_payload_corrupt      ), //i
    .io_ups_1_d_valid           (peripheral_bus_arbiter_core_io_ups_1_d_valid                   ), //o
    .io_ups_1_d_ready           (splited_mBus_to_peripheral_bus_down_bus_d_ready                ), //i
    .io_ups_1_d_payload_opcode  (peripheral_bus_arbiter_core_io_ups_1_d_payload_opcode[2:0]     ), //o
    .io_ups_1_d_payload_param   (peripheral_bus_arbiter_core_io_ups_1_d_payload_param[2:0]      ), //o
    .io_ups_1_d_payload_source  (peripheral_bus_arbiter_core_io_ups_1_d_payload_source[1:0]     ), //o
    .io_ups_1_d_payload_size    (peripheral_bus_arbiter_core_io_ups_1_d_payload_size[2:0]       ), //o
    .io_ups_1_d_payload_denied  (peripheral_bus_arbiter_core_io_ups_1_d_payload_denied          ), //o
    .io_ups_1_d_payload_data    (peripheral_bus_arbiter_core_io_ups_1_d_payload_data[31:0]      ), //o
    .io_ups_1_d_payload_corrupt (peripheral_bus_arbiter_core_io_ups_1_d_payload_corrupt         ), //o
    .io_down_a_valid            (peripheral_bus_arbiter_core_io_down_a_valid                    ), //o
    .io_down_a_ready            (peripheral_bus_bus_a_ready                                     ), //i
    .io_down_a_payload_opcode   (peripheral_bus_arbiter_core_io_down_a_payload_opcode[2:0]      ), //o
    .io_down_a_payload_param    (peripheral_bus_arbiter_core_io_down_a_payload_param[2:0]       ), //o
    .io_down_a_payload_source   (peripheral_bus_arbiter_core_io_down_a_payload_source[2:0]      ), //o
    .io_down_a_payload_address  (peripheral_bus_arbiter_core_io_down_a_payload_address[31:0]    ), //o
    .io_down_a_payload_size     (peripheral_bus_arbiter_core_io_down_a_payload_size[2:0]        ), //o
    .io_down_a_payload_mask     (peripheral_bus_arbiter_core_io_down_a_payload_mask[3:0]        ), //o
    .io_down_a_payload_data     (peripheral_bus_arbiter_core_io_down_a_payload_data[31:0]       ), //o
    .io_down_a_payload_corrupt  (peripheral_bus_arbiter_core_io_down_a_payload_corrupt          ), //o
    .io_down_d_valid            (peripheral_bus_bus_d_valid                                     ), //i
    .io_down_d_ready            (peripheral_bus_arbiter_core_io_down_d_ready                    ), //o
    .io_down_d_payload_opcode   (peripheral_bus_bus_d_payload_opcode[2:0]                       ), //i
    .io_down_d_payload_param    (peripheral_bus_bus_d_payload_param[2:0]                        ), //i
    .io_down_d_payload_source   (peripheral_bus_bus_d_payload_source[2:0]                       ), //i
    .io_down_d_payload_size     (peripheral_bus_bus_d_payload_size[2:0]                         ), //i
    .io_down_d_payload_denied   (peripheral_bus_bus_d_payload_denied                            ), //i
    .io_down_d_payload_data     (peripheral_bus_bus_d_payload_data[31:0]                        ), //i
    .io_down_d_payload_corrupt  (peripheral_bus_bus_d_payload_corrupt                           ), //i
    .litex_clk                  (litex_clk                                                      ), //i
    .litex_reset                (litex_reset                                                    )  //i
  );
  Axi4Bridge mem_toAxi4_logic_bridge (
    .io_up_a_valid              (mem_toAxi4_up_bus_a_valid                            ), //i
    .io_up_a_ready              (mem_toAxi4_logic_bridge_io_up_a_ready                ), //o
    .io_up_a_payload_opcode     (mem_toAxi4_up_bus_a_payload_opcode[2:0]              ), //i
    .io_up_a_payload_param      (mem_toAxi4_up_bus_a_payload_param[2:0]               ), //i
    .io_up_a_payload_source     (mem_toAxi4_up_bus_a_payload_source[1:0]              ), //i
    .io_up_a_payload_address    (mem_toAxi4_up_bus_a_payload_address[31:0]            ), //i
    .io_up_a_payload_size       (mem_toAxi4_up_bus_a_payload_size[2:0]                ), //i
    .io_up_a_payload_mask       (mem_toAxi4_up_bus_a_payload_mask[15:0]               ), //i
    .io_up_a_payload_data       (mem_toAxi4_up_bus_a_payload_data[127:0]              ), //i
    .io_up_a_payload_corrupt    (mem_toAxi4_up_bus_a_payload_corrupt                  ), //i
    .io_up_d_valid              (mem_toAxi4_logic_bridge_io_up_d_valid                ), //o
    .io_up_d_ready              (mem_toAxi4_up_bus_d_ready                            ), //i
    .io_up_d_payload_opcode     (mem_toAxi4_logic_bridge_io_up_d_payload_opcode[2:0]  ), //o
    .io_up_d_payload_param      (mem_toAxi4_logic_bridge_io_up_d_payload_param[2:0]   ), //o
    .io_up_d_payload_source     (mem_toAxi4_logic_bridge_io_up_d_payload_source[1:0]  ), //o
    .io_up_d_payload_size       (mem_toAxi4_logic_bridge_io_up_d_payload_size[2:0]    ), //o
    .io_up_d_payload_denied     (mem_toAxi4_logic_bridge_io_up_d_payload_denied       ), //o
    .io_up_d_payload_data       (mem_toAxi4_logic_bridge_io_up_d_payload_data[127:0]  ), //o
    .io_up_d_payload_corrupt    (mem_toAxi4_logic_bridge_io_up_d_payload_corrupt      ), //o
    .io_down_aw_valid           (mem_toAxi4_logic_bridge_io_down_aw_valid             ), //o
    .io_down_aw_ready           (mem_toAxi4_down_aw_ready                             ), //i
    .io_down_aw_payload_addr    (mem_toAxi4_logic_bridge_io_down_aw_payload_addr[31:0]), //o
    .io_down_aw_payload_id      (mem_toAxi4_logic_bridge_io_down_aw_payload_id[1:0]   ), //o
    .io_down_aw_payload_len     (mem_toAxi4_logic_bridge_io_down_aw_payload_len[7:0]  ), //o
    .io_down_aw_payload_size    (mem_toAxi4_logic_bridge_io_down_aw_payload_size[2:0] ), //o
    .io_down_aw_payload_burst   (mem_toAxi4_logic_bridge_io_down_aw_payload_burst[1:0]), //o
    .io_down_aw_payload_allStrb (mem_toAxi4_logic_bridge_io_down_aw_payload_allStrb   ), //o
    .io_down_w_valid            (mem_toAxi4_logic_bridge_io_down_w_valid              ), //o
    .io_down_w_ready            (mem_toAxi4_down_w_ready                              ), //i
    .io_down_w_payload_data     (mem_toAxi4_logic_bridge_io_down_w_payload_data[127:0]), //o
    .io_down_w_payload_strb     (mem_toAxi4_logic_bridge_io_down_w_payload_strb[15:0] ), //o
    .io_down_w_payload_last     (mem_toAxi4_logic_bridge_io_down_w_payload_last       ), //o
    .io_down_b_valid            (mem_toAxi4_down_b_valid                              ), //i
    .io_down_b_ready            (mem_toAxi4_logic_bridge_io_down_b_ready              ), //o
    .io_down_b_payload_id       (mem_toAxi4_down_b_payload_id[1:0]                    ), //i
    .io_down_b_payload_resp     (mem_toAxi4_down_b_payload_resp[1:0]                  ), //i
    .io_down_ar_valid           (mem_toAxi4_logic_bridge_io_down_ar_valid             ), //o
    .io_down_ar_ready           (mem_toAxi4_down_ar_ready                             ), //i
    .io_down_ar_payload_addr    (mem_toAxi4_logic_bridge_io_down_ar_payload_addr[31:0]), //o
    .io_down_ar_payload_id      (mem_toAxi4_logic_bridge_io_down_ar_payload_id[1:0]   ), //o
    .io_down_ar_payload_len     (mem_toAxi4_logic_bridge_io_down_ar_payload_len[7:0]  ), //o
    .io_down_ar_payload_size    (mem_toAxi4_logic_bridge_io_down_ar_payload_size[2:0] ), //o
    .io_down_ar_payload_burst   (mem_toAxi4_logic_bridge_io_down_ar_payload_burst[1:0]), //o
    .io_down_r_valid            (mem_toAxi4_down_r_valid                              ), //i
    .io_down_r_ready            (mem_toAxi4_logic_bridge_io_down_r_ready              ), //o
    .io_down_r_payload_data     (mem_toAxi4_down_r_payload_data[127:0]                ), //i
    .io_down_r_payload_id       (mem_toAxi4_down_r_payload_id[1:0]                    ), //i
    .io_down_r_payload_resp     (mem_toAxi4_down_r_payload_resp[1:0]                  ), //i
    .io_down_r_payload_last     (mem_toAxi4_down_r_payload_last                       ), //i
    .litex_clk                  (litex_clk                                            ), //i
    .cpuResetCtrl_reset         (cpuResetCtrl_reset                                   )  //i
  );
  Decoder splited_mBus_decoder_core (
    .io_up_a_valid                (splited_mBus_bus_a_valid                                    ), //i
    .io_up_a_ready                (splited_mBus_decoder_core_io_up_a_ready                     ), //o
    .io_up_a_payload_opcode       (splited_mBus_bus_a_payload_opcode[2:0]                      ), //i
    .io_up_a_payload_param        (splited_mBus_bus_a_payload_param[2:0]                       ), //i
    .io_up_a_payload_source       (splited_mBus_bus_a_payload_source[1:0]                      ), //i
    .io_up_a_payload_address      (splited_mBus_bus_a_payload_address[31:0]                    ), //i
    .io_up_a_payload_size         (splited_mBus_bus_a_payload_size[2:0]                        ), //i
    .io_up_a_payload_mask         (splited_mBus_bus_a_payload_mask[7:0]                        ), //i
    .io_up_a_payload_data         (splited_mBus_bus_a_payload_data[63:0]                       ), //i
    .io_up_a_payload_corrupt      (splited_mBus_bus_a_payload_corrupt                          ), //i
    .io_up_d_valid                (splited_mBus_decoder_core_io_up_d_valid                     ), //o
    .io_up_d_ready                (splited_mBus_bus_d_ready                                    ), //i
    .io_up_d_payload_opcode       (splited_mBus_decoder_core_io_up_d_payload_opcode[2:0]       ), //o
    .io_up_d_payload_param        (splited_mBus_decoder_core_io_up_d_payload_param[2:0]        ), //o
    .io_up_d_payload_source       (splited_mBus_decoder_core_io_up_d_payload_source[1:0]       ), //o
    .io_up_d_payload_size         (splited_mBus_decoder_core_io_up_d_payload_size[2:0]         ), //o
    .io_up_d_payload_denied       (splited_mBus_decoder_core_io_up_d_payload_denied            ), //o
    .io_up_d_payload_data         (splited_mBus_decoder_core_io_up_d_payload_data[63:0]        ), //o
    .io_up_d_payload_corrupt      (splited_mBus_decoder_core_io_up_d_payload_corrupt           ), //o
    .io_downs_0_a_valid           (splited_mBus_decoder_core_io_downs_0_a_valid                ), //o
    .io_downs_0_a_ready           (splited_mBus_to_mem_toAxi4_up_up_bus_a_ready                ), //i
    .io_downs_0_a_payload_opcode  (splited_mBus_decoder_core_io_downs_0_a_payload_opcode[2:0]  ), //o
    .io_downs_0_a_payload_param   (splited_mBus_decoder_core_io_downs_0_a_payload_param[2:0]   ), //o
    .io_downs_0_a_payload_source  (splited_mBus_decoder_core_io_downs_0_a_payload_source[1:0]  ), //o
    .io_downs_0_a_payload_address (splited_mBus_decoder_core_io_downs_0_a_payload_address[31:0]), //o
    .io_downs_0_a_payload_size    (splited_mBus_decoder_core_io_downs_0_a_payload_size[2:0]    ), //o
    .io_downs_0_a_payload_mask    (splited_mBus_decoder_core_io_downs_0_a_payload_mask[7:0]    ), //o
    .io_downs_0_a_payload_data    (splited_mBus_decoder_core_io_downs_0_a_payload_data[63:0]   ), //o
    .io_downs_0_a_payload_corrupt (splited_mBus_decoder_core_io_downs_0_a_payload_corrupt      ), //o
    .io_downs_0_d_valid           (splited_mBus_to_mem_toAxi4_up_up_bus_d_valid                ), //i
    .io_downs_0_d_ready           (splited_mBus_decoder_core_io_downs_0_d_ready                ), //o
    .io_downs_0_d_payload_opcode  (splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode[2:0]  ), //i
    .io_downs_0_d_payload_param   (splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_param[2:0]   ), //i
    .io_downs_0_d_payload_source  (splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_source[1:0]  ), //i
    .io_downs_0_d_payload_size    (splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_size[2:0]    ), //i
    .io_downs_0_d_payload_denied  (splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_denied       ), //i
    .io_downs_0_d_payload_data    (splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_data[63:0]   ), //i
    .io_downs_0_d_payload_corrupt (splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_corrupt      ), //i
    .io_downs_1_a_valid           (splited_mBus_decoder_core_io_downs_1_a_valid                ), //o
    .io_downs_1_a_ready           (splited_mBus_to_peripheral_bus_up_bus_a_ready               ), //i
    .io_downs_1_a_payload_opcode  (splited_mBus_decoder_core_io_downs_1_a_payload_opcode[2:0]  ), //o
    .io_downs_1_a_payload_param   (splited_mBus_decoder_core_io_downs_1_a_payload_param[2:0]   ), //o
    .io_downs_1_a_payload_source  (splited_mBus_decoder_core_io_downs_1_a_payload_source[1:0]  ), //o
    .io_downs_1_a_payload_address (splited_mBus_decoder_core_io_downs_1_a_payload_address[31:0]), //o
    .io_downs_1_a_payload_size    (splited_mBus_decoder_core_io_downs_1_a_payload_size[2:0]    ), //o
    .io_downs_1_a_payload_mask    (splited_mBus_decoder_core_io_downs_1_a_payload_mask[7:0]    ), //o
    .io_downs_1_a_payload_data    (splited_mBus_decoder_core_io_downs_1_a_payload_data[63:0]   ), //o
    .io_downs_1_a_payload_corrupt (splited_mBus_decoder_core_io_downs_1_a_payload_corrupt      ), //o
    .io_downs_1_d_valid           (splited_mBus_to_peripheral_bus_up_bus_d_valid               ), //i
    .io_downs_1_d_ready           (splited_mBus_decoder_core_io_downs_1_d_ready                ), //o
    .io_downs_1_d_payload_opcode  (splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode[2:0] ), //i
    .io_downs_1_d_payload_param   (splited_mBus_to_peripheral_bus_up_bus_d_payload_param[2:0]  ), //i
    .io_downs_1_d_payload_source  (splited_mBus_to_peripheral_bus_up_bus_d_payload_source[1:0] ), //i
    .io_downs_1_d_payload_size    (splited_mBus_to_peripheral_bus_up_bus_d_payload_size[2:0]   ), //i
    .io_downs_1_d_payload_denied  (splited_mBus_to_peripheral_bus_up_bus_d_payload_denied      ), //i
    .io_downs_1_d_payload_data    (splited_mBus_to_peripheral_bus_up_bus_d_payload_data[63:0]  ), //i
    .io_downs_1_d_payload_corrupt (splited_mBus_to_peripheral_bus_up_bus_d_payload_corrupt     ), //i
    .litex_clk                    (litex_clk                                                   ), //i
    .cpuResetCtrl_reset           (cpuResetCtrl_reset                                          )  //i
  );
  TilelinkClint peripheral_clint_thread_core (
    .io_bus_a_valid           (peripheral_clint_node_bus_a_valid                        ), //i
    .io_bus_a_ready           (peripheral_clint_thread_core_io_bus_a_ready              ), //o
    .io_bus_a_payload_opcode  (peripheral_clint_node_bus_a_payload_opcode[2:0]          ), //i
    .io_bus_a_payload_param   (peripheral_clint_node_bus_a_payload_param[2:0]           ), //i
    .io_bus_a_payload_source  (peripheral_clint_node_bus_a_payload_source[2:0]          ), //i
    .io_bus_a_payload_address (peripheral_clint_node_bus_a_payload_address[15:0]        ), //i
    .io_bus_a_payload_size    (peripheral_clint_node_bus_a_payload_size[2:0]            ), //i
    .io_bus_a_payload_mask    (peripheral_clint_node_bus_a_payload_mask[3:0]            ), //i
    .io_bus_a_payload_data    (peripheral_clint_node_bus_a_payload_data[31:0]           ), //i
    .io_bus_a_payload_corrupt (peripheral_clint_node_bus_a_payload_corrupt              ), //i
    .io_bus_d_valid           (peripheral_clint_thread_core_io_bus_d_valid              ), //o
    .io_bus_d_ready           (peripheral_clint_node_bus_d_ready                        ), //i
    .io_bus_d_payload_opcode  (peripheral_clint_thread_core_io_bus_d_payload_opcode[2:0]), //o
    .io_bus_d_payload_param   (peripheral_clint_thread_core_io_bus_d_payload_param[2:0] ), //o
    .io_bus_d_payload_source  (peripheral_clint_thread_core_io_bus_d_payload_source[2:0]), //o
    .io_bus_d_payload_size    (peripheral_clint_thread_core_io_bus_d_payload_size[2:0]  ), //o
    .io_bus_d_payload_denied  (peripheral_clint_thread_core_io_bus_d_payload_denied     ), //o
    .io_bus_d_payload_data    (peripheral_clint_thread_core_io_bus_d_payload_data[31:0] ), //o
    .io_bus_d_payload_corrupt (peripheral_clint_thread_core_io_bus_d_payload_corrupt    ), //o
    .io_timerInterrupt        (peripheral_clint_thread_core_io_timerInterrupt           ), //o
    .io_softwareInterrupt     (peripheral_clint_thread_core_io_softwareInterrupt        ), //o
    .io_time                  (peripheral_clint_thread_core_io_time[63:0]               ), //o
    .io_stop                  (peripheral_clint_thread_core_io_stop                     ), //i
    .litex_clk                (litex_clk                                                ), //i
    .litex_reset              (litex_reset                                              )  //i
  );
  TilelinkPlic peripheral_plic_thread_logic (
    .io_bus_a_valid           (peripheral_plic_node_bus_a_valid                         ), //i
    .io_bus_a_ready           (peripheral_plic_thread_logic_io_bus_a_ready              ), //o
    .io_bus_a_payload_opcode  (peripheral_plic_node_bus_a_payload_opcode[2:0]           ), //i
    .io_bus_a_payload_param   (peripheral_plic_node_bus_a_payload_param[2:0]            ), //i
    .io_bus_a_payload_source  (peripheral_plic_node_bus_a_payload_source[2:0]           ), //i
    .io_bus_a_payload_address (peripheral_plic_node_bus_a_payload_address[21:0]         ), //i
    .io_bus_a_payload_size    (peripheral_plic_node_bus_a_payload_size[1:0]             ), //i
    .io_bus_a_payload_mask    (peripheral_plic_node_bus_a_payload_mask[3:0]             ), //i
    .io_bus_a_payload_data    (peripheral_plic_node_bus_a_payload_data[31:0]            ), //i
    .io_bus_a_payload_corrupt (peripheral_plic_node_bus_a_payload_corrupt               ), //i
    .io_bus_d_valid           (peripheral_plic_thread_logic_io_bus_d_valid              ), //o
    .io_bus_d_ready           (peripheral_plic_node_bus_d_ready                         ), //i
    .io_bus_d_payload_opcode  (peripheral_plic_thread_logic_io_bus_d_payload_opcode[2:0]), //o
    .io_bus_d_payload_param   (peripheral_plic_thread_logic_io_bus_d_payload_param[2:0] ), //o
    .io_bus_d_payload_source  (peripheral_plic_thread_logic_io_bus_d_payload_source[2:0]), //o
    .io_bus_d_payload_size    (peripheral_plic_thread_logic_io_bus_d_payload_size[1:0]  ), //o
    .io_bus_d_payload_denied  (peripheral_plic_thread_logic_io_bus_d_payload_denied     ), //o
    .io_bus_d_payload_data    (peripheral_plic_thread_logic_io_bus_d_payload_data[31:0] ), //o
    .io_bus_d_payload_corrupt (peripheral_plic_thread_logic_io_bus_d_payload_corrupt    ), //o
    .io_sources               (peripheral_plic_thread_logic_io_sources[30:0]            ), //i
    .io_targets               (peripheral_plic_thread_logic_io_targets[1:0]             ), //o
    .litex_clk                (litex_clk                                                ), //i
    .litex_reset              (litex_reset                                              )  //i
  );
  AxiLite4Bridge peripheral_toAxiLite4_logic_bridge (
    .io_up_a_valid           (peripheral_toAxiLite4_up_bus_a_valid                            ), //i
    .io_up_a_ready           (peripheral_toAxiLite4_logic_bridge_io_up_a_ready                ), //o
    .io_up_a_payload_opcode  (peripheral_toAxiLite4_up_bus_a_payload_opcode[2:0]              ), //i
    .io_up_a_payload_param   (peripheral_toAxiLite4_up_bus_a_payload_param[2:0]               ), //i
    .io_up_a_payload_source  (peripheral_toAxiLite4_up_bus_a_payload_source[2:0]              ), //i
    .io_up_a_payload_address (peripheral_toAxiLite4_up_bus_a_payload_address[31:0]            ), //i
    .io_up_a_payload_size    (peripheral_toAxiLite4_up_bus_a_payload_size[2:0]                ), //i
    .io_up_a_payload_mask    (peripheral_toAxiLite4_up_bus_a_payload_mask[3:0]                ), //i
    .io_up_a_payload_data    (peripheral_toAxiLite4_up_bus_a_payload_data[31:0]               ), //i
    .io_up_a_payload_corrupt (peripheral_toAxiLite4_up_bus_a_payload_corrupt                  ), //i
    .io_up_d_valid           (peripheral_toAxiLite4_logic_bridge_io_up_d_valid                ), //o
    .io_up_d_ready           (peripheral_toAxiLite4_up_bus_d_ready                            ), //i
    .io_up_d_payload_opcode  (peripheral_toAxiLite4_logic_bridge_io_up_d_payload_opcode[2:0]  ), //o
    .io_up_d_payload_param   (peripheral_toAxiLite4_logic_bridge_io_up_d_payload_param[2:0]   ), //o
    .io_up_d_payload_source  (peripheral_toAxiLite4_logic_bridge_io_up_d_payload_source[2:0]  ), //o
    .io_up_d_payload_size    (peripheral_toAxiLite4_logic_bridge_io_up_d_payload_size[2:0]    ), //o
    .io_up_d_payload_denied  (peripheral_toAxiLite4_logic_bridge_io_up_d_payload_denied       ), //o
    .io_up_d_payload_data    (peripheral_toAxiLite4_logic_bridge_io_up_d_payload_data[31:0]   ), //o
    .io_up_d_payload_corrupt (peripheral_toAxiLite4_logic_bridge_io_up_d_payload_corrupt      ), //o
    .io_down_aw_valid        (peripheral_toAxiLite4_logic_bridge_io_down_aw_valid             ), //o
    .io_down_aw_ready        (peripheral_toAxiLite4_down_aw_ready                             ), //i
    .io_down_aw_payload_addr (peripheral_toAxiLite4_logic_bridge_io_down_aw_payload_addr[31:0]), //o
    .io_down_aw_payload_prot (peripheral_toAxiLite4_logic_bridge_io_down_aw_payload_prot[2:0] ), //o
    .io_down_w_valid         (peripheral_toAxiLite4_logic_bridge_io_down_w_valid              ), //o
    .io_down_w_ready         (peripheral_toAxiLite4_down_w_ready                              ), //i
    .io_down_w_payload_data  (peripheral_toAxiLite4_logic_bridge_io_down_w_payload_data[31:0] ), //o
    .io_down_w_payload_strb  (peripheral_toAxiLite4_logic_bridge_io_down_w_payload_strb[3:0]  ), //o
    .io_down_b_valid         (peripheral_toAxiLite4_down_b_valid                              ), //i
    .io_down_b_ready         (peripheral_toAxiLite4_logic_bridge_io_down_b_ready              ), //o
    .io_down_b_payload_resp  (peripheral_toAxiLite4_down_b_payload_resp[1:0]                  ), //i
    .io_down_ar_valid        (peripheral_toAxiLite4_logic_bridge_io_down_ar_valid             ), //o
    .io_down_ar_ready        (peripheral_toAxiLite4_down_ar_ready                             ), //i
    .io_down_ar_payload_addr (peripheral_toAxiLite4_logic_bridge_io_down_ar_payload_addr[31:0]), //o
    .io_down_ar_payload_prot (peripheral_toAxiLite4_logic_bridge_io_down_ar_payload_prot[2:0] ), //o
    .io_down_r_valid         (peripheral_toAxiLite4_down_r_valid                              ), //i
    .io_down_r_ready         (peripheral_toAxiLite4_logic_bridge_io_down_r_ready              ), //o
    .io_down_r_payload_data  (peripheral_toAxiLite4_down_r_payload_data[31:0]                 ), //i
    .io_down_r_payload_resp  (peripheral_toAxiLite4_down_r_payload_resp[1:0]                  ), //i
    .litex_clk               (litex_clk                                                       ), //i
    .litex_reset             (litex_reset                                                     )  //i
  );
  WidthAdapter splited_mBus_to_mem_toAxi4_up_widthAdapter (
    .io_up_a_valid             (splited_mBus_to_mem_toAxi4_up_up_bus_a_valid                              ), //i
    .io_up_a_ready             (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_a_ready                  ), //o
    .io_up_a_payload_opcode    (splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode[2:0]                ), //i
    .io_up_a_payload_param     (splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_param[2:0]                 ), //i
    .io_up_a_payload_source    (splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_source[1:0]                ), //i
    .io_up_a_payload_address   (splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_address[31:0]              ), //i
    .io_up_a_payload_size      (splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_size[2:0]                  ), //i
    .io_up_a_payload_mask      (splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_mask[7:0]                  ), //i
    .io_up_a_payload_data      (splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_data[63:0]                 ), //i
    .io_up_a_payload_corrupt   (splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_corrupt                    ), //i
    .io_up_d_valid             (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_valid                  ), //o
    .io_up_d_ready             (splited_mBus_to_mem_toAxi4_up_up_bus_d_ready                              ), //i
    .io_up_d_payload_opcode    (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_opcode[2:0]    ), //o
    .io_up_d_payload_param     (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_param[2:0]     ), //o
    .io_up_d_payload_source    (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_source[1:0]    ), //o
    .io_up_d_payload_size      (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_size[2:0]      ), //o
    .io_up_d_payload_denied    (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_denied         ), //o
    .io_up_d_payload_data      (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_data[63:0]     ), //o
    .io_up_d_payload_corrupt   (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_corrupt        ), //o
    .io_down_a_valid           (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_valid                ), //o
    .io_down_a_ready           (splited_mBus_to_mem_toAxi4_up_down_bus_a_ready                            ), //i
    .io_down_a_payload_opcode  (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_opcode[2:0]  ), //o
    .io_down_a_payload_param   (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_param[2:0]   ), //o
    .io_down_a_payload_source  (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_source[1:0]  ), //o
    .io_down_a_payload_address (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_address[31:0]), //o
    .io_down_a_payload_size    (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_size[2:0]    ), //o
    .io_down_a_payload_mask    (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_mask[15:0]   ), //o
    .io_down_a_payload_data    (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_data[127:0]  ), //o
    .io_down_a_payload_corrupt (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_corrupt      ), //o
    .io_down_d_valid           (splited_mBus_to_mem_toAxi4_up_down_bus_d_valid                            ), //i
    .io_down_d_ready           (splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_d_ready                ), //o
    .io_down_d_payload_opcode  (splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode[2:0]              ), //i
    .io_down_d_payload_param   (splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_param[2:0]               ), //i
    .io_down_d_payload_source  (splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_source[1:0]              ), //i
    .io_down_d_payload_size    (splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_size[2:0]                ), //i
    .io_down_d_payload_denied  (splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_denied                   ), //i
    .io_down_d_payload_data    (splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_data[127:0]              ), //i
    .io_down_d_payload_corrupt (splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_corrupt                  ), //i
    .litex_clk                 (litex_clk                                                                 ), //i
    .cpuResetCtrl_reset        (cpuResetCtrl_reset                                                        )  //i
  );
  WidthAdapter_1 splited_mBus_to_peripheral_bus_widthAdapter (
    .io_up_a_valid             (splited_mBus_to_peripheral_bus_up_bus_a_valid                              ), //i
    .io_up_a_ready             (splited_mBus_to_peripheral_bus_widthAdapter_io_up_a_ready                  ), //o
    .io_up_a_payload_opcode    (splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode[2:0]                ), //i
    .io_up_a_payload_param     (splited_mBus_to_peripheral_bus_up_bus_a_payload_param[2:0]                 ), //i
    .io_up_a_payload_source    (splited_mBus_to_peripheral_bus_up_bus_a_payload_source[1:0]                ), //i
    .io_up_a_payload_address   (splited_mBus_to_peripheral_bus_up_bus_a_payload_address[31:0]              ), //i
    .io_up_a_payload_size      (splited_mBus_to_peripheral_bus_up_bus_a_payload_size[2:0]                  ), //i
    .io_up_a_payload_mask      (splited_mBus_to_peripheral_bus_up_bus_a_payload_mask[7:0]                  ), //i
    .io_up_a_payload_data      (splited_mBus_to_peripheral_bus_up_bus_a_payload_data[63:0]                 ), //i
    .io_up_a_payload_corrupt   (splited_mBus_to_peripheral_bus_up_bus_a_payload_corrupt                    ), //i
    .io_up_d_valid             (splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_valid                  ), //o
    .io_up_d_ready             (splited_mBus_to_peripheral_bus_up_bus_d_ready                              ), //i
    .io_up_d_payload_opcode    (splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_opcode[2:0]    ), //o
    .io_up_d_payload_param     (splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_param[2:0]     ), //o
    .io_up_d_payload_source    (splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_source[1:0]    ), //o
    .io_up_d_payload_size      (splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_size[2:0]      ), //o
    .io_up_d_payload_denied    (splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_denied         ), //o
    .io_up_d_payload_data      (splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_data[63:0]     ), //o
    .io_up_d_payload_corrupt   (splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_corrupt        ), //o
    .io_down_a_valid           (splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_valid                ), //o
    .io_down_a_ready           (splited_mBus_to_peripheral_bus_down_bus_a_ready                            ), //i
    .io_down_a_payload_opcode  (splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_opcode[2:0]  ), //o
    .io_down_a_payload_param   (splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_param[2:0]   ), //o
    .io_down_a_payload_source  (splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_source[1:0]  ), //o
    .io_down_a_payload_address (splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_address[31:0]), //o
    .io_down_a_payload_size    (splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_size[2:0]    ), //o
    .io_down_a_payload_mask    (splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_mask[3:0]    ), //o
    .io_down_a_payload_data    (splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_data[31:0]   ), //o
    .io_down_a_payload_corrupt (splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_corrupt      ), //o
    .io_down_d_valid           (splited_mBus_to_peripheral_bus_down_bus_d_valid                            ), //i
    .io_down_d_ready           (splited_mBus_to_peripheral_bus_widthAdapter_io_down_d_ready                ), //o
    .io_down_d_payload_opcode  (splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode[2:0]              ), //i
    .io_down_d_payload_param   (splited_mBus_to_peripheral_bus_down_bus_d_payload_param[2:0]               ), //i
    .io_down_d_payload_source  (splited_mBus_to_peripheral_bus_down_bus_d_payload_source[1:0]              ), //i
    .io_down_d_payload_size    (splited_mBus_to_peripheral_bus_down_bus_d_payload_size[2:0]                ), //i
    .io_down_d_payload_denied  (splited_mBus_to_peripheral_bus_down_bus_d_payload_denied                   ), //i
    .io_down_d_payload_data    (splited_mBus_to_peripheral_bus_down_bus_d_payload_data[31:0]               ), //i
    .io_down_d_payload_corrupt (splited_mBus_to_peripheral_bus_down_bus_d_payload_corrupt                  ), //i
    .litex_clk                 (litex_clk                                                                  ), //i
    .litex_reset               (litex_reset                                                                )  //i
  );
  Decoder_1 peripheral_bus_decoder_core (
    .io_up_a_valid                (peripheral_bus_bus_a_halfPipe_valid                                    ), //i
    .io_up_a_ready                (peripheral_bus_decoder_core_io_up_a_ready                              ), //o
    .io_up_a_payload_opcode       (peripheral_bus_bus_a_halfPipe_payload_opcode[2:0]                      ), //i
    .io_up_a_payload_param        (peripheral_bus_bus_a_halfPipe_payload_param[2:0]                       ), //i
    .io_up_a_payload_source       (peripheral_bus_bus_a_halfPipe_payload_source[2:0]                      ), //i
    .io_up_a_payload_address      (peripheral_bus_bus_a_halfPipe_payload_address[31:0]                    ), //i
    .io_up_a_payload_size         (peripheral_bus_bus_a_halfPipe_payload_size[2:0]                        ), //i
    .io_up_a_payload_mask         (peripheral_bus_bus_a_halfPipe_payload_mask[3:0]                        ), //i
    .io_up_a_payload_data         (peripheral_bus_bus_a_halfPipe_payload_data[31:0]                       ), //i
    .io_up_a_payload_corrupt      (peripheral_bus_bus_a_halfPipe_payload_corrupt                          ), //i
    .io_up_d_valid                (peripheral_bus_decoder_core_io_up_d_valid                              ), //o
    .io_up_d_ready                (peripheral_bus_decoder_core_io_up_d_ready                              ), //i
    .io_up_d_payload_opcode       (peripheral_bus_decoder_core_io_up_d_payload_opcode[2:0]                ), //o
    .io_up_d_payload_param        (peripheral_bus_decoder_core_io_up_d_payload_param[2:0]                 ), //o
    .io_up_d_payload_source       (peripheral_bus_decoder_core_io_up_d_payload_source[2:0]                ), //o
    .io_up_d_payload_size         (peripheral_bus_decoder_core_io_up_d_payload_size[2:0]                  ), //o
    .io_up_d_payload_denied       (peripheral_bus_decoder_core_io_up_d_payload_denied                     ), //o
    .io_up_d_payload_data         (peripheral_bus_decoder_core_io_up_d_payload_data[31:0]                 ), //o
    .io_up_d_payload_corrupt      (peripheral_bus_decoder_core_io_up_d_payload_corrupt                    ), //o
    .io_downs_0_a_valid           (peripheral_bus_decoder_core_io_downs_0_a_valid                         ), //o
    .io_downs_0_a_ready           (peripheral_bus_to_peripheral_clint_node_up_bus_a_ready                 ), //i
    .io_downs_0_a_payload_opcode  (peripheral_bus_decoder_core_io_downs_0_a_payload_opcode[2:0]           ), //o
    .io_downs_0_a_payload_param   (peripheral_bus_decoder_core_io_downs_0_a_payload_param[2:0]            ), //o
    .io_downs_0_a_payload_source  (peripheral_bus_decoder_core_io_downs_0_a_payload_source[2:0]           ), //o
    .io_downs_0_a_payload_address (peripheral_bus_decoder_core_io_downs_0_a_payload_address[15:0]         ), //o
    .io_downs_0_a_payload_size    (peripheral_bus_decoder_core_io_downs_0_a_payload_size[2:0]             ), //o
    .io_downs_0_a_payload_mask    (peripheral_bus_decoder_core_io_downs_0_a_payload_mask[3:0]             ), //o
    .io_downs_0_a_payload_data    (peripheral_bus_decoder_core_io_downs_0_a_payload_data[31:0]            ), //o
    .io_downs_0_a_payload_corrupt (peripheral_bus_decoder_core_io_downs_0_a_payload_corrupt               ), //o
    .io_downs_0_d_valid           (peripheral_bus_to_peripheral_clint_node_up_bus_d_valid                 ), //i
    .io_downs_0_d_ready           (peripheral_bus_decoder_core_io_downs_0_d_ready                         ), //o
    .io_downs_0_d_payload_opcode  (peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode[2:0]   ), //i
    .io_downs_0_d_payload_param   (peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_param[2:0]    ), //i
    .io_downs_0_d_payload_source  (peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_source[2:0]   ), //i
    .io_downs_0_d_payload_size    (peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_size[2:0]     ), //i
    .io_downs_0_d_payload_denied  (peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_denied        ), //i
    .io_downs_0_d_payload_data    (peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_data[31:0]    ), //i
    .io_downs_0_d_payload_corrupt (peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_corrupt       ), //i
    .io_downs_1_a_valid           (peripheral_bus_decoder_core_io_downs_1_a_valid                         ), //o
    .io_downs_1_a_ready           (peripheral_bus_to_peripheral_plic_node_up_bus_a_ready                  ), //i
    .io_downs_1_a_payload_opcode  (peripheral_bus_decoder_core_io_downs_1_a_payload_opcode[2:0]           ), //o
    .io_downs_1_a_payload_param   (peripheral_bus_decoder_core_io_downs_1_a_payload_param[2:0]            ), //o
    .io_downs_1_a_payload_source  (peripheral_bus_decoder_core_io_downs_1_a_payload_source[2:0]           ), //o
    .io_downs_1_a_payload_address (peripheral_bus_decoder_core_io_downs_1_a_payload_address[21:0]         ), //o
    .io_downs_1_a_payload_size    (peripheral_bus_decoder_core_io_downs_1_a_payload_size[1:0]             ), //o
    .io_downs_1_a_payload_mask    (peripheral_bus_decoder_core_io_downs_1_a_payload_mask[3:0]             ), //o
    .io_downs_1_a_payload_data    (peripheral_bus_decoder_core_io_downs_1_a_payload_data[31:0]            ), //o
    .io_downs_1_a_payload_corrupt (peripheral_bus_decoder_core_io_downs_1_a_payload_corrupt               ), //o
    .io_downs_1_d_valid           (peripheral_bus_to_peripheral_plic_node_up_bus_d_valid                  ), //i
    .io_downs_1_d_ready           (peripheral_bus_decoder_core_io_downs_1_d_ready                         ), //o
    .io_downs_1_d_payload_opcode  (peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode[2:0]    ), //i
    .io_downs_1_d_payload_param   (peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_param[2:0]     ), //i
    .io_downs_1_d_payload_source  (peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_source[2:0]    ), //i
    .io_downs_1_d_payload_size    (peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_size[1:0]      ), //i
    .io_downs_1_d_payload_denied  (peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_denied         ), //i
    .io_downs_1_d_payload_data    (peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_data[31:0]     ), //i
    .io_downs_1_d_payload_corrupt (peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_corrupt        ), //i
    .io_downs_2_a_valid           (peripheral_bus_decoder_core_io_downs_2_a_valid                         ), //o
    .io_downs_2_a_ready           (peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_ready              ), //i
    .io_downs_2_a_payload_opcode  (peripheral_bus_decoder_core_io_downs_2_a_payload_opcode[2:0]           ), //o
    .io_downs_2_a_payload_param   (peripheral_bus_decoder_core_io_downs_2_a_payload_param[2:0]            ), //o
    .io_downs_2_a_payload_source  (peripheral_bus_decoder_core_io_downs_2_a_payload_source[2:0]           ), //o
    .io_downs_2_a_payload_address (peripheral_bus_decoder_core_io_downs_2_a_payload_address[31:0]         ), //o
    .io_downs_2_a_payload_size    (peripheral_bus_decoder_core_io_downs_2_a_payload_size[2:0]             ), //o
    .io_downs_2_a_payload_mask    (peripheral_bus_decoder_core_io_downs_2_a_payload_mask[3:0]             ), //o
    .io_downs_2_a_payload_data    (peripheral_bus_decoder_core_io_downs_2_a_payload_data[31:0]            ), //o
    .io_downs_2_a_payload_corrupt (peripheral_bus_decoder_core_io_downs_2_a_payload_corrupt               ), //o
    .io_downs_2_d_valid           (peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_valid              ), //i
    .io_downs_2_d_ready           (peripheral_bus_decoder_core_io_downs_2_d_ready                         ), //o
    .io_downs_2_d_payload_opcode  (peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode[2:0]), //i
    .io_downs_2_d_payload_param   (peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_param[2:0] ), //i
    .io_downs_2_d_payload_source  (peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_source[2:0]), //i
    .io_downs_2_d_payload_size    (peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_size[2:0]  ), //i
    .io_downs_2_d_payload_denied  (peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_denied     ), //i
    .io_downs_2_d_payload_data    (peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_data[31:0] ), //i
    .io_downs_2_d_payload_corrupt (peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_corrupt    ), //i
    .litex_clk                    (litex_clk                                                              ), //i
    .litex_reset                  (litex_reset                                                            )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(vexiis_0_dBus_bus_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_dBus_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_dBus_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_dBus_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_dBus_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_dBus_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_dBus_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_bus_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_dBus_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_dBus_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_dBus_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_dBus_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_dBus_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_dBus_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_noDecoder_toDown_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_dBus_noDecoder_toDown_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_dBus_noDecoder_toDown_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_dBus_noDecoder_toDown_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_dBus_noDecoder_toDown_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_dBus_noDecoder_toDown_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_dBus_noDecoder_toDown_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_noDecoder_toDown_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_dBus_noDecoder_toDown_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_dBus_noDecoder_toDown_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_dBus_noDecoder_toDown_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_dBus_noDecoder_toDown_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_dBus_noDecoder_toDown_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_dBus_noDecoder_toDown_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_bus_a_halfPipe_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_dBus_bus_a_halfPipe_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_dBus_bus_a_halfPipe_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_dBus_bus_a_halfPipe_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_dBus_bus_a_halfPipe_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_dBus_bus_a_halfPipe_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_dBus_bus_a_halfPipe_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_bus_a_rData_opcode)
      A_PUT_FULL_DATA : vexiis_0_dBus_bus_a_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_dBus_bus_a_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_dBus_bus_a_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_dBus_bus_a_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_dBus_bus_a_rData_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_dBus_bus_a_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode)
      D_ACCESS_ACK : vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_noDecoder_toDown_d_rData_opcode)
      D_ACCESS_ACK : vexiis_0_dBus_noDecoder_toDown_d_rData_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_dBus_noDecoder_toDown_d_rData_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_dBus_noDecoder_toDown_d_rData_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_dBus_noDecoder_toDown_d_rData_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_dBus_noDecoder_toDown_d_rData_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_dBus_noDecoder_toDown_d_rData_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_bus_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_iBus_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_iBus_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_iBus_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_iBus_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_iBus_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_iBus_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_bus_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_iBus_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_iBus_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_iBus_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_iBus_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_iBus_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_iBus_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_noDecoder_toDown_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_iBus_noDecoder_toDown_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_iBus_noDecoder_toDown_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_iBus_noDecoder_toDown_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_iBus_noDecoder_toDown_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_iBus_noDecoder_toDown_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_iBus_noDecoder_toDown_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_noDecoder_toDown_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_iBus_noDecoder_toDown_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_iBus_noDecoder_toDown_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_iBus_noDecoder_toDown_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_iBus_noDecoder_toDown_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_iBus_noDecoder_toDown_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_iBus_noDecoder_toDown_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_bus_a_halfPipe_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_iBus_bus_a_halfPipe_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_iBus_bus_a_halfPipe_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_iBus_bus_a_halfPipe_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_iBus_bus_a_halfPipe_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_iBus_bus_a_halfPipe_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_iBus_bus_a_halfPipe_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_bus_a_rData_opcode)
      A_PUT_FULL_DATA : vexiis_0_iBus_bus_a_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_iBus_bus_a_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_iBus_bus_a_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_iBus_bus_a_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_iBus_bus_a_rData_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_iBus_bus_a_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_bus_a_halfPipe_rData_opcode)
      A_PUT_FULL_DATA : vexiis_0_iBus_bus_a_halfPipe_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_iBus_bus_a_halfPipe_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_iBus_bus_a_halfPipe_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_iBus_bus_a_halfPipe_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_iBus_bus_a_halfPipe_rData_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_iBus_bus_a_halfPipe_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_noDecoder_connection_payload_opcode)
      D_ACCESS_ACK : vexiis_0_iBus_noDecoder_connection_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_iBus_noDecoder_connection_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_iBus_noDecoder_connection_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_iBus_noDecoder_connection_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_iBus_noDecoder_connection_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_iBus_noDecoder_connection_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_noDecoder_toDown_d_rData_opcode)
      D_ACCESS_ACK : vexiis_0_iBus_noDecoder_toDown_d_rData_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_iBus_noDecoder_toDown_d_rData_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_iBus_noDecoder_toDown_d_rData_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_iBus_noDecoder_toDown_d_rData_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_iBus_noDecoder_toDown_d_rData_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_iBus_noDecoder_toDown_d_rData_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_bus_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_lsuL1Bus_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_lsuL1Bus_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_lsuL1Bus_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_lsuL1Bus_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_lsuL1Bus_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_lsuL1Bus_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_bus_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_lsuL1Bus_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_lsuL1Bus_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_lsuL1Bus_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_lsuL1Bus_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_lsuL1Bus_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_lsuL1Bus_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_bus_a_rData_opcode)
      A_PUT_FULL_DATA : vexiis_0_lsuL1Bus_bus_a_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_lsuL1Bus_bus_a_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_lsuL1Bus_bus_a_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_lsuL1Bus_bus_a_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_lsuL1Bus_bus_a_rData_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_lsuL1Bus_bus_a_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode)
      A_PUT_FULL_DATA : _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode)
      A_PUT_FULL_DATA : vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode)
      D_ACCESS_ACK : vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode)
      D_ACCESS_ACK : vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ioBus_bus_a_payload_opcode)
      A_PUT_FULL_DATA : ioBus_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ioBus_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ioBus_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ioBus_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ioBus_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ioBus_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ioBus_bus_d_payload_opcode)
      D_ACCESS_ACK : ioBus_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ioBus_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ioBus_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ioBus_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ioBus_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ioBus_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode)
      A_PUT_FULL_DATA : vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ioBus_bus_d_combStage_payload_opcode)
      D_ACCESS_ACK : ioBus_bus_d_combStage_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ioBus_bus_d_combStage_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ioBus_bus_d_combStage_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ioBus_bus_d_combStage_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ioBus_bus_d_combStage_payload_opcode_string = "RELEASE_ACK    ";
      default : ioBus_bus_d_combStage_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ioBus_noDecoder_toDown_a_payload_opcode)
      A_PUT_FULL_DATA : ioBus_noDecoder_toDown_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ioBus_noDecoder_toDown_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ioBus_noDecoder_toDown_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ioBus_noDecoder_toDown_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ioBus_noDecoder_toDown_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ioBus_noDecoder_toDown_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ioBus_noDecoder_toDown_d_payload_opcode)
      D_ACCESS_ACK : ioBus_noDecoder_toDown_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ioBus_noDecoder_toDown_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ioBus_noDecoder_toDown_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ioBus_noDecoder_toDown_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ioBus_noDecoder_toDown_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ioBus_noDecoder_toDown_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_bus_a_payload_opcode)
      A_PUT_FULL_DATA : splited_mBus_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : splited_mBus_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : splited_mBus_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : splited_mBus_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : splited_mBus_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : splited_mBus_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_bus_d_payload_opcode)
      D_ACCESS_ACK : splited_mBus_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : splited_mBus_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : splited_mBus_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : splited_mBus_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : splited_mBus_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : splited_mBus_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_bus_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_bus_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_bus_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_bus_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_bus_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_bus_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_bus_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_bus_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_bus_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_bus_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_bus_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_bus_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ioBus_to_peripheral_bus_down_bus_a_payload_opcode)
      A_PUT_FULL_DATA : ioBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ioBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ioBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ioBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ioBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ioBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ioBus_to_peripheral_bus_down_bus_d_payload_opcode)
      D_ACCESS_ACK : ioBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ioBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ioBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ioBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ioBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ioBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode)
      A_PUT_FULL_DATA : splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode)
      D_ACCESS_ACK : splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(mem_toAxi4_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : mem_toAxi4_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : mem_toAxi4_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : mem_toAxi4_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : mem_toAxi4_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : mem_toAxi4_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : mem_toAxi4_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(mem_toAxi4_up_bus_d_payload_opcode)
      D_ACCESS_ACK : mem_toAxi4_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : mem_toAxi4_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : mem_toAxi4_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : mem_toAxi4_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : mem_toAxi4_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : mem_toAxi4_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode)
      A_PUT_FULL_DATA : splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode)
      D_ACCESS_ACK : splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode)
      D_ACCESS_ACK : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_clint_node_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_clint_node_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_clint_node_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_clint_node_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_clint_node_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_clint_node_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_clint_node_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_clint_node_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_clint_node_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_clint_node_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_clint_node_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_clint_node_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_clint_node_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_clint_node_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_plic_node_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_plic_node_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_plic_node_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_plic_node_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_plic_node_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_plic_node_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_plic_node_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_plic_node_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_plic_node_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_plic_node_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_plic_node_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_plic_node_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_plic_node_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_plic_node_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_toAxiLite4_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_toAxiLite4_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_toAxiLite4_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_toAxiLite4_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_toAxiLite4_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_toAxiLite4_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_toAxiLite4_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_toAxiLite4_up_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_toAxiLite4_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_toAxiLite4_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_toAxiLite4_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_toAxiLite4_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_toAxiLite4_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_toAxiLite4_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ioBus_to_peripheral_bus_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : ioBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ioBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ioBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ioBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ioBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ioBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ioBus_to_peripheral_bus_up_bus_d_payload_opcode)
      D_ACCESS_ACK : ioBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ioBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ioBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ioBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ioBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ioBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode)
      D_ACCESS_ACK : splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode)
      D_ACCESS_ACK : splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode)
      A_PUT_FULL_DATA : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode)
      D_ACCESS_ACK : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_bus_a_halfPipe_payload_opcode)
      A_PUT_FULL_DATA : peripheral_bus_bus_a_halfPipe_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_bus_bus_a_halfPipe_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_bus_bus_a_halfPipe_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_bus_bus_a_halfPipe_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_bus_bus_a_halfPipe_payload_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_bus_bus_a_halfPipe_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(peripheral_bus_bus_a_rData_opcode)
      A_PUT_FULL_DATA : peripheral_bus_bus_a_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : peripheral_bus_bus_a_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : peripheral_bus_bus_a_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : peripheral_bus_bus_a_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : peripheral_bus_bus_a_rData_opcode_string = "ACQUIRE_PERM    ";
      default : peripheral_bus_bus_a_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_halfPipe_payload_opcode)
      D_ACCESS_ACK : io_up_d_halfPipe_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_halfPipe_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_halfPipe_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_halfPipe_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_halfPipe_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_halfPipe_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_rData_opcode)
      D_ACCESS_ACK : io_up_d_rData_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_rData_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_rData_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_rData_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_rData_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_rData_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign peripheral_externalInterrupts_toPlic_1_node_flag = peripheral_externalInterrupts_port[1];
  assign peripheral_externalInterrupts_toPlic_2_node_flag = peripheral_externalInterrupts_port[2];
  assign peripheral_externalInterrupts_toPlic_3_node_flag = peripheral_externalInterrupts_port[3];
  assign peripheral_externalInterrupts_toPlic_4_node_flag = peripheral_externalInterrupts_port[4];
  assign peripheral_externalInterrupts_toPlic_5_node_flag = peripheral_externalInterrupts_port[5];
  assign peripheral_externalInterrupts_toPlic_6_node_flag = peripheral_externalInterrupts_port[6];
  assign peripheral_externalInterrupts_toPlic_7_node_flag = peripheral_externalInterrupts_port[7];
  assign peripheral_externalInterrupts_toPlic_8_node_flag = peripheral_externalInterrupts_port[8];
  assign peripheral_externalInterrupts_toPlic_9_node_flag = peripheral_externalInterrupts_port[9];
  assign peripheral_externalInterrupts_toPlic_10_node_flag = peripheral_externalInterrupts_port[10];
  assign peripheral_externalInterrupts_toPlic_11_node_flag = peripheral_externalInterrupts_port[11];
  assign peripheral_externalInterrupts_toPlic_12_node_flag = peripheral_externalInterrupts_port[12];
  assign peripheral_externalInterrupts_toPlic_13_node_flag = peripheral_externalInterrupts_port[13];
  assign peripheral_externalInterrupts_toPlic_14_node_flag = peripheral_externalInterrupts_port[14];
  assign peripheral_externalInterrupts_toPlic_15_node_flag = peripheral_externalInterrupts_port[15];
  assign peripheral_externalInterrupts_toPlic_16_node_flag = peripheral_externalInterrupts_port[16];
  assign peripheral_externalInterrupts_toPlic_17_node_flag = peripheral_externalInterrupts_port[17];
  assign peripheral_externalInterrupts_toPlic_18_node_flag = peripheral_externalInterrupts_port[18];
  assign peripheral_externalInterrupts_toPlic_19_node_flag = peripheral_externalInterrupts_port[19];
  assign peripheral_externalInterrupts_toPlic_20_node_flag = peripheral_externalInterrupts_port[20];
  assign peripheral_externalInterrupts_toPlic_21_node_flag = peripheral_externalInterrupts_port[21];
  assign peripheral_externalInterrupts_toPlic_22_node_flag = peripheral_externalInterrupts_port[22];
  assign peripheral_externalInterrupts_toPlic_23_node_flag = peripheral_externalInterrupts_port[23];
  assign peripheral_externalInterrupts_toPlic_24_node_flag = peripheral_externalInterrupts_port[24];
  assign peripheral_externalInterrupts_toPlic_25_node_flag = peripheral_externalInterrupts_port[25];
  assign peripheral_externalInterrupts_toPlic_26_node_flag = peripheral_externalInterrupts_port[26];
  assign peripheral_externalInterrupts_toPlic_27_node_flag = peripheral_externalInterrupts_port[27];
  assign peripheral_externalInterrupts_toPlic_28_node_flag = peripheral_externalInterrupts_port[28];
  assign peripheral_externalInterrupts_toPlic_29_node_flag = peripheral_externalInterrupts_port[29];
  assign peripheral_externalInterrupts_toPlic_30_node_flag = peripheral_externalInterrupts_port[30];
  assign peripheral_externalInterrupts_toPlic_31_node_flag = peripheral_externalInterrupts_port[31];
  assign vexiis_0_priv_rdtime = _zz_vexiis_0_priv_rdtime;
  assign cpuResetCtrl_fiber_aggregator_reset = (|cpuResetCtrl_fiber_aggregator_asyncBuffers_0_io_dataOut);
  assign cpuResetCtrl_fiber_holder_reset = ((cpuResetCtrl_fiber_holder_counter != 7'h40) ^ 1'b0);
  assign when_CrossClock_l341 = (cpuResetCtrl_fiber_holder_reset == 1'b1);
  assign cpuResetCtrl_reset = cpuResetCtrl_fiber_buffer_io_dataOut;
  assign vexiis_0_priv_mti_thread_gateways_0_flag = peripheral_clint_thread_core_io_timerInterrupt[0];
  assign vexiis_0_priv_mti_flag = (|vexiis_0_priv_mti_thread_gateways_0_flag);
  assign vexiis_0_priv_msi_thread_gateways_0_flag = peripheral_clint_thread_core_io_softwareInterrupt[0];
  assign vexiis_0_priv_msi_flag = (|vexiis_0_priv_msi_thread_gateways_0_flag);
  assign vexiis_0_priv_mei_thread_gateways_0_flag = peripheral_plic_to_vexiis_0_priv_mei_flag;
  assign vexiis_0_priv_mei_flag = (|vexiis_0_priv_mei_thread_gateways_0_flag);
  assign vexiis_0_priv_sei_thread_gateways_0_flag = peripheral_plic_to_vexiis_0_priv_sei_flag;
  assign vexiis_0_priv_sei_flag = (|vexiis_0_priv_sei_thread_gateways_0_flag);
  assign vexiis_0_dBus_bus_a_halfPipe_fire = (vexiis_0_dBus_bus_a_halfPipe_valid && vexiis_0_dBus_bus_a_halfPipe_ready);
  assign vexiis_0_dBus_bus_a_ready = (! vexiis_0_dBus_bus_a_rValid);
  assign vexiis_0_dBus_bus_a_halfPipe_valid = vexiis_0_dBus_bus_a_rValid;
  assign vexiis_0_dBus_bus_a_halfPipe_payload_opcode = vexiis_0_dBus_bus_a_rData_opcode;
  assign vexiis_0_dBus_bus_a_halfPipe_payload_param = vexiis_0_dBus_bus_a_rData_param;
  assign vexiis_0_dBus_bus_a_halfPipe_payload_address = vexiis_0_dBus_bus_a_rData_address;
  assign vexiis_0_dBus_bus_a_halfPipe_payload_size = vexiis_0_dBus_bus_a_rData_size;
  assign vexiis_0_dBus_bus_a_halfPipe_payload_mask = vexiis_0_dBus_bus_a_rData_mask;
  assign vexiis_0_dBus_bus_a_halfPipe_payload_data = vexiis_0_dBus_bus_a_rData_data;
  assign vexiis_0_dBus_bus_a_halfPipe_payload_corrupt = vexiis_0_dBus_bus_a_rData_corrupt;
  assign vexiis_0_dBus_noDecoder_toDown_a_valid = vexiis_0_dBus_bus_a_halfPipe_valid;
  assign vexiis_0_dBus_bus_a_halfPipe_ready = vexiis_0_dBus_noDecoder_toDown_a_ready;
  assign vexiis_0_dBus_noDecoder_toDown_a_payload_opcode = vexiis_0_dBus_bus_a_halfPipe_payload_opcode;
  assign vexiis_0_dBus_noDecoder_toDown_a_payload_param = vexiis_0_dBus_bus_a_halfPipe_payload_param;
  assign vexiis_0_dBus_noDecoder_toDown_a_payload_address = vexiis_0_dBus_bus_a_halfPipe_payload_address;
  assign vexiis_0_dBus_noDecoder_toDown_a_payload_size = vexiis_0_dBus_bus_a_halfPipe_payload_size;
  assign vexiis_0_dBus_noDecoder_toDown_a_payload_mask = vexiis_0_dBus_bus_a_halfPipe_payload_mask;
  assign vexiis_0_dBus_noDecoder_toDown_a_payload_data = vexiis_0_dBus_bus_a_halfPipe_payload_data;
  assign vexiis_0_dBus_noDecoder_toDown_a_payload_corrupt = vexiis_0_dBus_bus_a_halfPipe_payload_corrupt;
  always @(*) begin
    vexiis_0_dBus_noDecoder_toDown_d_ready = vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_ready;
    if(when_Stream_l399) begin
      vexiis_0_dBus_noDecoder_toDown_d_ready = 1'b1;
    end
  end

  assign when_Stream_l399 = (! vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_valid);
  assign vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_valid = vexiis_0_dBus_noDecoder_toDown_d_rValid;
  assign vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode = vexiis_0_dBus_noDecoder_toDown_d_rData_opcode;
  assign vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_param = vexiis_0_dBus_noDecoder_toDown_d_rData_param;
  assign vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_size = vexiis_0_dBus_noDecoder_toDown_d_rData_size;
  assign vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_denied = vexiis_0_dBus_noDecoder_toDown_d_rData_denied;
  assign vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_data = vexiis_0_dBus_noDecoder_toDown_d_rData_data;
  assign vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_corrupt = vexiis_0_dBus_noDecoder_toDown_d_rData_corrupt;
  assign vexiis_0_dBus_bus_d_valid = vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_valid;
  assign vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_ready = vexiis_0_dBus_bus_d_ready;
  assign vexiis_0_dBus_bus_d_payload_opcode = vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_opcode;
  assign vexiis_0_dBus_bus_d_payload_param = vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_param;
  assign vexiis_0_dBus_bus_d_payload_size = vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_size;
  assign vexiis_0_dBus_bus_d_payload_denied = vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_denied;
  assign vexiis_0_dBus_bus_d_payload_data = vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_data;
  assign vexiis_0_dBus_bus_d_payload_corrupt = vexiis_0_dBus_noDecoder_toDown_d_m2sPipe_payload_corrupt;
  assign vexiis_0_iBus_bus_a_halfPipe_fire = (vexiis_0_iBus_bus_a_halfPipe_valid && vexiis_0_iBus_bus_a_halfPipe_ready);
  assign vexiis_0_iBus_bus_a_ready = (! vexiis_0_iBus_bus_a_rValid);
  assign vexiis_0_iBus_bus_a_halfPipe_valid = vexiis_0_iBus_bus_a_rValid;
  assign vexiis_0_iBus_bus_a_halfPipe_payload_opcode = vexiis_0_iBus_bus_a_rData_opcode;
  assign vexiis_0_iBus_bus_a_halfPipe_payload_param = vexiis_0_iBus_bus_a_rData_param;
  assign vexiis_0_iBus_bus_a_halfPipe_payload_address = vexiis_0_iBus_bus_a_rData_address;
  assign vexiis_0_iBus_bus_a_halfPipe_payload_size = vexiis_0_iBus_bus_a_rData_size;
  assign vexiis_0_iBus_bus_a_halfPipe_halfPipe_fire = (vexiis_0_iBus_bus_a_halfPipe_halfPipe_valid && vexiis_0_iBus_bus_a_halfPipe_halfPipe_ready);
  assign vexiis_0_iBus_bus_a_halfPipe_ready = (! vexiis_0_iBus_bus_a_halfPipe_rValid);
  assign vexiis_0_iBus_bus_a_halfPipe_halfPipe_valid = vexiis_0_iBus_bus_a_halfPipe_rValid;
  assign vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode = vexiis_0_iBus_bus_a_halfPipe_rData_opcode;
  assign vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_param = vexiis_0_iBus_bus_a_halfPipe_rData_param;
  assign vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_address = vexiis_0_iBus_bus_a_halfPipe_rData_address;
  assign vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_size = vexiis_0_iBus_bus_a_halfPipe_rData_size;
  assign vexiis_0_iBus_noDecoder_toDown_a_valid = vexiis_0_iBus_bus_a_halfPipe_halfPipe_valid;
  assign vexiis_0_iBus_bus_a_halfPipe_halfPipe_ready = vexiis_0_iBus_noDecoder_toDown_a_ready;
  assign vexiis_0_iBus_noDecoder_toDown_a_payload_opcode = vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_opcode;
  assign vexiis_0_iBus_noDecoder_toDown_a_payload_param = vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_param;
  assign vexiis_0_iBus_noDecoder_toDown_a_payload_address = vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_address;
  assign vexiis_0_iBus_noDecoder_toDown_a_payload_size = vexiis_0_iBus_bus_a_halfPipe_halfPipe_payload_size;
  always @(*) begin
    vexiis_0_iBus_noDecoder_toDown_d_ready = vexiis_0_iBus_noDecoder_connection_ready;
    if(when_Stream_l399_1) begin
      vexiis_0_iBus_noDecoder_toDown_d_ready = 1'b1;
    end
  end

  assign when_Stream_l399_1 = (! vexiis_0_iBus_noDecoder_connection_valid);
  assign vexiis_0_iBus_noDecoder_connection_valid = vexiis_0_iBus_noDecoder_toDown_d_rValid;
  assign vexiis_0_iBus_noDecoder_connection_payload_opcode = vexiis_0_iBus_noDecoder_toDown_d_rData_opcode;
  assign vexiis_0_iBus_noDecoder_connection_payload_param = vexiis_0_iBus_noDecoder_toDown_d_rData_param;
  assign vexiis_0_iBus_noDecoder_connection_payload_size = vexiis_0_iBus_noDecoder_toDown_d_rData_size;
  assign vexiis_0_iBus_noDecoder_connection_payload_denied = vexiis_0_iBus_noDecoder_toDown_d_rData_denied;
  assign vexiis_0_iBus_noDecoder_connection_payload_data = vexiis_0_iBus_noDecoder_toDown_d_rData_data;
  assign vexiis_0_iBus_noDecoder_connection_payload_corrupt = vexiis_0_iBus_noDecoder_toDown_d_rData_corrupt;
  assign vexiis_0_iBus_bus_d_valid = vexiis_0_iBus_noDecoder_connection_valid;
  assign vexiis_0_iBus_noDecoder_connection_ready = vexiis_0_iBus_bus_d_ready;
  assign vexiis_0_iBus_bus_d_payload_opcode = vexiis_0_iBus_noDecoder_connection_payload_opcode;
  assign vexiis_0_iBus_bus_d_payload_param = vexiis_0_iBus_noDecoder_connection_payload_param;
  assign vexiis_0_iBus_bus_d_payload_size = vexiis_0_iBus_noDecoder_connection_payload_size;
  assign vexiis_0_iBus_bus_d_payload_denied = vexiis_0_iBus_noDecoder_connection_payload_denied;
  assign vexiis_0_iBus_bus_d_payload_data = vexiis_0_iBus_noDecoder_connection_payload_data;
  assign vexiis_0_iBus_bus_d_payload_corrupt = vexiis_0_iBus_noDecoder_connection_payload_corrupt;
  assign vexiis_0_lsuL1Bus_bus_a_ready = vexiis_0_lsuL1Bus_bus_a_rValidN;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_valid = (vexiis_0_lsuL1Bus_bus_a_valid || (! vexiis_0_lsuL1Bus_bus_a_rValidN));
  assign _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode = (vexiis_0_lsuL1Bus_bus_a_rValidN ? vexiis_0_lsuL1Bus_bus_a_payload_opcode : vexiis_0_lsuL1Bus_bus_a_rData_opcode);
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode = _zz_vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_param = (vexiis_0_lsuL1Bus_bus_a_rValidN ? vexiis_0_lsuL1Bus_bus_a_payload_param : vexiis_0_lsuL1Bus_bus_a_rData_param);
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_source = (vexiis_0_lsuL1Bus_bus_a_rValidN ? vexiis_0_lsuL1Bus_bus_a_payload_source : vexiis_0_lsuL1Bus_bus_a_rData_source);
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_address = (vexiis_0_lsuL1Bus_bus_a_rValidN ? vexiis_0_lsuL1Bus_bus_a_payload_address : vexiis_0_lsuL1Bus_bus_a_rData_address);
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_size = (vexiis_0_lsuL1Bus_bus_a_rValidN ? vexiis_0_lsuL1Bus_bus_a_payload_size : vexiis_0_lsuL1Bus_bus_a_rData_size);
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_mask = (vexiis_0_lsuL1Bus_bus_a_rValidN ? vexiis_0_lsuL1Bus_bus_a_payload_mask : vexiis_0_lsuL1Bus_bus_a_rData_mask);
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_data = (vexiis_0_lsuL1Bus_bus_a_rValidN ? vexiis_0_lsuL1Bus_bus_a_payload_data : vexiis_0_lsuL1Bus_bus_a_rData_data);
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_corrupt = (vexiis_0_lsuL1Bus_bus_a_rValidN ? vexiis_0_lsuL1Bus_bus_a_payload_corrupt : vexiis_0_lsuL1Bus_bus_a_rData_corrupt);
  always @(*) begin
    vexiis_0_lsuL1Bus_bus_a_s2mPipe_ready = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_ready;
    if(when_Stream_l399_2) begin
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l399_2 = (! vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_valid);
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_valid = vexiis_0_lsuL1Bus_bus_a_s2mPipe_rValid;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode = vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_param = vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_param;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_source = vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_source;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_address = vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_address;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_size = vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_size;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_mask = vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_mask;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_data = vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_data;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_corrupt = vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_corrupt;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_valid = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_valid;
  assign vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_ready = vexiis_0_lsuL1Bus_noDecoder_toDown_a_ready;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_opcode;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_param = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_param;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_source = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_source;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_address = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_address;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_size = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_size;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_mask = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_mask;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_data = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_data;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_corrupt = vexiis_0_lsuL1Bus_bus_a_s2mPipe_m2sPipe_payload_corrupt;
  always @(*) begin
    vexiis_0_lsuL1Bus_noDecoder_toDown_d_ready = vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_ready;
    if(when_Stream_l399_3) begin
      vexiis_0_lsuL1Bus_noDecoder_toDown_d_ready = 1'b1;
    end
  end

  assign when_Stream_l399_3 = (! vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_valid);
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_valid = vexiis_0_lsuL1Bus_noDecoder_toDown_d_rValid;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode = vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_param = vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_param;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_source = vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_source;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_size = vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_size;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_denied = vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_denied;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_data = vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_data;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_corrupt = vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_corrupt;
  assign vexiis_0_lsuL1Bus_bus_d_valid = vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_valid;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_ready = vexiis_0_lsuL1Bus_bus_d_ready;
  assign vexiis_0_lsuL1Bus_bus_d_payload_opcode = vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_opcode;
  assign vexiis_0_lsuL1Bus_bus_d_payload_param = vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_param;
  assign vexiis_0_lsuL1Bus_bus_d_payload_source = vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_source;
  assign vexiis_0_lsuL1Bus_bus_d_payload_size = vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_size;
  assign vexiis_0_lsuL1Bus_bus_d_payload_denied = vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_denied;
  assign vexiis_0_lsuL1Bus_bus_d_payload_data = vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_data;
  assign vexiis_0_lsuL1Bus_bus_d_payload_corrupt = vexiis_0_lsuL1Bus_noDecoder_toDown_d_m2sPipe_payload_corrupt;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_fire = (vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_valid && vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_ready);
  assign vexiis_0_dBus_to_ioBus_down_bus_a_ready = (! vexiis_0_dBus_to_ioBus_down_bus_a_rValid);
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_valid = vexiis_0_dBus_to_ioBus_down_bus_a_rValid;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode = vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_param = vexiis_0_dBus_to_ioBus_down_bus_a_rData_param;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_address = vexiis_0_dBus_to_ioBus_down_bus_a_rData_address;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_size = vexiis_0_dBus_to_ioBus_down_bus_a_rData_size;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_mask = vexiis_0_dBus_to_ioBus_down_bus_a_rData_mask;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_data = vexiis_0_dBus_to_ioBus_down_bus_a_rData_data;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_corrupt = vexiis_0_dBus_to_ioBus_down_bus_a_rData_corrupt;
  assign ioBus_bus_a_valid = vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_valid;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_ready = ioBus_bus_a_ready;
  assign ioBus_bus_a_payload_opcode = vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_opcode;
  assign ioBus_bus_a_payload_param = vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_param;
  assign ioBus_bus_a_payload_address = vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_address;
  assign ioBus_bus_a_payload_size = vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_size;
  assign ioBus_bus_a_payload_mask = vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_mask;
  assign ioBus_bus_a_payload_data = vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_data;
  assign ioBus_bus_a_payload_corrupt = vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_payload_corrupt;
  assign ioBus_bus_d_combStage_valid = ioBus_bus_d_valid;
  assign ioBus_bus_d_ready = ioBus_bus_d_combStage_ready;
  assign ioBus_bus_d_combStage_payload_opcode = ioBus_bus_d_payload_opcode;
  assign ioBus_bus_d_combStage_payload_param = ioBus_bus_d_payload_param;
  assign ioBus_bus_d_combStage_payload_size = ioBus_bus_d_payload_size;
  assign ioBus_bus_d_combStage_payload_denied = ioBus_bus_d_payload_denied;
  assign ioBus_bus_d_combStage_payload_data = ioBus_bus_d_payload_data;
  assign ioBus_bus_d_combStage_payload_corrupt = ioBus_bus_d_payload_corrupt;
  assign vexiis_0_dBus_to_ioBus_down_bus_d_valid = ioBus_bus_d_combStage_valid;
  assign ioBus_bus_d_combStage_ready = vexiis_0_dBus_to_ioBus_down_bus_d_ready;
  assign vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode = ioBus_bus_d_combStage_payload_opcode;
  assign vexiis_0_dBus_to_ioBus_down_bus_d_payload_param = ioBus_bus_d_combStage_payload_param;
  assign vexiis_0_dBus_to_ioBus_down_bus_d_payload_size = ioBus_bus_d_combStage_payload_size;
  assign vexiis_0_dBus_to_ioBus_down_bus_d_payload_denied = ioBus_bus_d_combStage_payload_denied;
  assign vexiis_0_dBus_to_ioBus_down_bus_d_payload_data = ioBus_bus_d_combStage_payload_data;
  assign vexiis_0_dBus_to_ioBus_down_bus_d_payload_corrupt = ioBus_bus_d_combStage_payload_corrupt;
  assign ioBus_noDecoder_toDown_a_valid = ioBus_bus_a_valid;
  assign ioBus_bus_a_ready = ioBus_noDecoder_toDown_a_ready;
  assign ioBus_noDecoder_toDown_a_payload_opcode = ioBus_bus_a_payload_opcode;
  assign ioBus_noDecoder_toDown_a_payload_param = ioBus_bus_a_payload_param;
  assign ioBus_noDecoder_toDown_a_payload_address = ioBus_bus_a_payload_address;
  assign ioBus_noDecoder_toDown_a_payload_size = ioBus_bus_a_payload_size;
  assign ioBus_noDecoder_toDown_a_payload_mask = ioBus_bus_a_payload_mask;
  assign ioBus_noDecoder_toDown_a_payload_data = ioBus_bus_a_payload_data;
  assign ioBus_noDecoder_toDown_a_payload_corrupt = ioBus_bus_a_payload_corrupt;
  assign ioBus_bus_d_valid = ioBus_noDecoder_toDown_d_valid;
  assign ioBus_noDecoder_toDown_d_ready = ioBus_bus_d_ready;
  assign ioBus_bus_d_payload_opcode = ioBus_noDecoder_toDown_d_payload_opcode;
  assign ioBus_bus_d_payload_param = ioBus_noDecoder_toDown_d_payload_param;
  assign ioBus_bus_d_payload_size = ioBus_noDecoder_toDown_d_payload_size;
  assign ioBus_bus_d_payload_denied = ioBus_noDecoder_toDown_d_payload_denied;
  assign ioBus_bus_d_payload_data = ioBus_noDecoder_toDown_d_payload_data;
  assign ioBus_bus_d_payload_corrupt = ioBus_noDecoder_toDown_d_payload_corrupt;
  assign vexiis_0_iBus_bus_a_valid = vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_valid;
  assign vexiis_0_iBus_bus_a_payload_opcode = vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_opcode;
  assign vexiis_0_iBus_bus_a_payload_param = vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_param;
  assign vexiis_0_iBus_bus_a_payload_address = vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_address;
  assign vexiis_0_iBus_bus_a_payload_size = vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_a_payload_size;
  assign vexiis_0_iBus_bus_d_ready = vexiis_0_logic_core_FetchL1TileLinkPlugin_logic_down_d_ready;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_a_ready = splited_mBus_arbiter_core_io_ups_0_a_ready;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_d_valid = splited_mBus_arbiter_core_io_ups_0_d_valid;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode = splited_mBus_arbiter_core_io_ups_0_d_payload_opcode;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_param = splited_mBus_arbiter_core_io_ups_0_d_payload_param;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_size = splited_mBus_arbiter_core_io_ups_0_d_payload_size;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_denied = splited_mBus_arbiter_core_io_ups_0_d_payload_denied;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_data = splited_mBus_arbiter_core_io_ups_0_d_payload_data;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_corrupt = splited_mBus_arbiter_core_io_ups_0_d_payload_corrupt;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_ready = splited_mBus_arbiter_core_io_ups_1_a_ready;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_valid = splited_mBus_arbiter_core_io_ups_1_d_valid;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode = splited_mBus_arbiter_core_io_ups_1_d_payload_opcode;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_param = splited_mBus_arbiter_core_io_ups_1_d_payload_param;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_source = splited_mBus_arbiter_core_io_ups_1_d_payload_source;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_size = splited_mBus_arbiter_core_io_ups_1_d_payload_size;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_denied = splited_mBus_arbiter_core_io_ups_1_d_payload_denied;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_data = splited_mBus_arbiter_core_io_ups_1_d_payload_data;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_corrupt = splited_mBus_arbiter_core_io_ups_1_d_payload_corrupt;
  assign splited_mBus_bus_a_valid = splited_mBus_arbiter_core_io_down_a_valid;
  assign splited_mBus_bus_a_payload_opcode = splited_mBus_arbiter_core_io_down_a_payload_opcode;
  assign splited_mBus_bus_a_payload_param = splited_mBus_arbiter_core_io_down_a_payload_param;
  assign splited_mBus_bus_a_payload_source = splited_mBus_arbiter_core_io_down_a_payload_source;
  assign splited_mBus_bus_a_payload_address = splited_mBus_arbiter_core_io_down_a_payload_address;
  assign splited_mBus_bus_a_payload_size = splited_mBus_arbiter_core_io_down_a_payload_size;
  assign splited_mBus_bus_a_payload_mask = splited_mBus_arbiter_core_io_down_a_payload_mask;
  assign splited_mBus_bus_a_payload_data = splited_mBus_arbiter_core_io_down_a_payload_data;
  assign splited_mBus_bus_a_payload_corrupt = splited_mBus_arbiter_core_io_down_a_payload_corrupt;
  assign splited_mBus_bus_d_ready = splited_mBus_arbiter_core_io_down_d_ready;
  assign ioBus_to_peripheral_bus_down_bus_a_ready = peripheral_bus_arbiter_core_io_ups_0_a_ready;
  assign ioBus_to_peripheral_bus_down_bus_d_valid = peripheral_bus_arbiter_core_io_ups_0_d_valid;
  assign ioBus_to_peripheral_bus_down_bus_d_payload_opcode = peripheral_bus_arbiter_core_io_ups_0_d_payload_opcode;
  assign ioBus_to_peripheral_bus_down_bus_d_payload_param = peripheral_bus_arbiter_core_io_ups_0_d_payload_param;
  assign ioBus_to_peripheral_bus_down_bus_d_payload_size = peripheral_bus_arbiter_core_io_ups_0_d_payload_size;
  assign ioBus_to_peripheral_bus_down_bus_d_payload_denied = peripheral_bus_arbiter_core_io_ups_0_d_payload_denied;
  assign ioBus_to_peripheral_bus_down_bus_d_payload_data = peripheral_bus_arbiter_core_io_ups_0_d_payload_data;
  assign ioBus_to_peripheral_bus_down_bus_d_payload_corrupt = peripheral_bus_arbiter_core_io_ups_0_d_payload_corrupt;
  assign splited_mBus_to_peripheral_bus_down_bus_a_ready = peripheral_bus_arbiter_core_io_ups_1_a_ready;
  assign splited_mBus_to_peripheral_bus_down_bus_d_valid = peripheral_bus_arbiter_core_io_ups_1_d_valid;
  assign splited_mBus_to_peripheral_bus_down_bus_d_payload_opcode = peripheral_bus_arbiter_core_io_ups_1_d_payload_opcode;
  assign splited_mBus_to_peripheral_bus_down_bus_d_payload_param = peripheral_bus_arbiter_core_io_ups_1_d_payload_param;
  assign splited_mBus_to_peripheral_bus_down_bus_d_payload_source = peripheral_bus_arbiter_core_io_ups_1_d_payload_source;
  assign splited_mBus_to_peripheral_bus_down_bus_d_payload_size = peripheral_bus_arbiter_core_io_ups_1_d_payload_size;
  assign splited_mBus_to_peripheral_bus_down_bus_d_payload_denied = peripheral_bus_arbiter_core_io_ups_1_d_payload_denied;
  assign splited_mBus_to_peripheral_bus_down_bus_d_payload_data = peripheral_bus_arbiter_core_io_ups_1_d_payload_data;
  assign splited_mBus_to_peripheral_bus_down_bus_d_payload_corrupt = peripheral_bus_arbiter_core_io_ups_1_d_payload_corrupt;
  assign peripheral_bus_bus_a_valid = peripheral_bus_arbiter_core_io_down_a_valid;
  assign peripheral_bus_bus_a_payload_opcode = peripheral_bus_arbiter_core_io_down_a_payload_opcode;
  assign peripheral_bus_bus_a_payload_param = peripheral_bus_arbiter_core_io_down_a_payload_param;
  assign peripheral_bus_bus_a_payload_source = peripheral_bus_arbiter_core_io_down_a_payload_source;
  assign peripheral_bus_bus_a_payload_address = peripheral_bus_arbiter_core_io_down_a_payload_address;
  assign peripheral_bus_bus_a_payload_size = peripheral_bus_arbiter_core_io_down_a_payload_size;
  assign peripheral_bus_bus_a_payload_mask = peripheral_bus_arbiter_core_io_down_a_payload_mask;
  assign peripheral_bus_bus_a_payload_data = peripheral_bus_arbiter_core_io_down_a_payload_data;
  assign peripheral_bus_bus_a_payload_corrupt = peripheral_bus_arbiter_core_io_down_a_payload_corrupt;
  assign peripheral_bus_bus_d_ready = peripheral_bus_arbiter_core_io_down_d_ready;
  assign vexiis_0_dBus_to_ioBus_up_bus_a_valid = vexiis_0_dBus_noDecoder_toDown_a_valid;
  assign vexiis_0_dBus_noDecoder_toDown_a_ready = vexiis_0_dBus_to_ioBus_up_bus_a_ready;
  assign vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode = vexiis_0_dBus_noDecoder_toDown_a_payload_opcode;
  assign vexiis_0_dBus_to_ioBus_up_bus_a_payload_param = vexiis_0_dBus_noDecoder_toDown_a_payload_param;
  assign vexiis_0_dBus_to_ioBus_up_bus_a_payload_mask = vexiis_0_dBus_noDecoder_toDown_a_payload_mask;
  assign vexiis_0_dBus_to_ioBus_up_bus_a_payload_data = vexiis_0_dBus_noDecoder_toDown_a_payload_data;
  assign vexiis_0_dBus_to_ioBus_up_bus_a_payload_corrupt = vexiis_0_dBus_noDecoder_toDown_a_payload_corrupt;
  assign vexiis_0_dBus_noDecoder_toDown_d_valid = vexiis_0_dBus_to_ioBus_up_bus_d_valid;
  assign vexiis_0_dBus_to_ioBus_up_bus_d_ready = vexiis_0_dBus_noDecoder_toDown_d_ready;
  assign vexiis_0_dBus_noDecoder_toDown_d_payload_opcode = vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode;
  assign vexiis_0_dBus_noDecoder_toDown_d_payload_param = vexiis_0_dBus_to_ioBus_up_bus_d_payload_param;
  assign vexiis_0_dBus_noDecoder_toDown_d_payload_denied = vexiis_0_dBus_to_ioBus_up_bus_d_payload_denied;
  assign vexiis_0_dBus_noDecoder_toDown_d_payload_data = vexiis_0_dBus_to_ioBus_up_bus_d_payload_data;
  assign vexiis_0_dBus_noDecoder_toDown_d_payload_corrupt = vexiis_0_dBus_to_ioBus_up_bus_d_payload_corrupt;
  assign vexiis_0_dBus_to_ioBus_up_bus_a_payload_size = vexiis_0_dBus_noDecoder_toDown_a_payload_size;
  assign vexiis_0_dBus_noDecoder_toDown_d_payload_size = vexiis_0_dBus_to_ioBus_up_bus_d_payload_size;
  assign vexiis_0_dBus_to_ioBus_up_bus_a_payload_address = vexiis_0_dBus_noDecoder_toDown_a_payload_address;
  assign vexiis_0_lsuL1Bus_bus_a_valid = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_valid;
  assign vexiis_0_lsuL1Bus_bus_a_payload_opcode = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_opcode;
  assign vexiis_0_lsuL1Bus_bus_a_payload_param = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_param;
  assign vexiis_0_lsuL1Bus_bus_a_payload_source = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_source;
  assign vexiis_0_lsuL1Bus_bus_a_payload_address = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_address;
  assign vexiis_0_lsuL1Bus_bus_a_payload_size = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_size;
  assign vexiis_0_lsuL1Bus_bus_a_payload_mask = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_mask;
  assign vexiis_0_lsuL1Bus_bus_a_payload_data = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_data;
  assign vexiis_0_lsuL1Bus_bus_a_payload_corrupt = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_a_payload_corrupt;
  assign vexiis_0_lsuL1Bus_bus_d_ready = vexiis_0_logic_core_LsuL1TileLinkPlugin_logic_down_d_ready;
  assign mem_toAxi4_up_bus_a_valid = splited_mBus_to_mem_toAxi4_up_down_bus_a_valid;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_ready = mem_toAxi4_up_bus_a_ready;
  assign mem_toAxi4_up_bus_a_payload_opcode = splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode;
  assign mem_toAxi4_up_bus_a_payload_param = splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_param;
  assign mem_toAxi4_up_bus_a_payload_source = splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_source;
  assign mem_toAxi4_up_bus_a_payload_address = splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_address;
  assign mem_toAxi4_up_bus_a_payload_size = splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_size;
  assign mem_toAxi4_up_bus_a_payload_mask = splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_mask;
  assign mem_toAxi4_up_bus_a_payload_data = splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_data;
  assign mem_toAxi4_up_bus_a_payload_corrupt = splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_corrupt;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_d_valid = mem_toAxi4_up_bus_d_valid;
  assign mem_toAxi4_up_bus_d_ready = splited_mBus_to_mem_toAxi4_up_down_bus_d_ready;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_opcode = mem_toAxi4_up_bus_d_payload_opcode;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_param = mem_toAxi4_up_bus_d_payload_param;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_source = mem_toAxi4_up_bus_d_payload_source;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_size = mem_toAxi4_up_bus_d_payload_size;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_denied = mem_toAxi4_up_bus_d_payload_denied;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_data = mem_toAxi4_up_bus_d_payload_data;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_d_payload_corrupt = mem_toAxi4_up_bus_d_payload_corrupt;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_a_valid = vexiis_0_iBus_noDecoder_toDown_a_valid;
  assign vexiis_0_iBus_noDecoder_toDown_a_ready = vexiis_0_iBus_to_splited_mBus_up_bus_a_ready;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode = vexiis_0_iBus_noDecoder_toDown_a_payload_opcode;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_param = vexiis_0_iBus_noDecoder_toDown_a_payload_param;
  assign vexiis_0_iBus_noDecoder_toDown_d_valid = vexiis_0_iBus_to_splited_mBus_up_bus_d_valid;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_d_ready = vexiis_0_iBus_noDecoder_toDown_d_ready;
  assign vexiis_0_iBus_noDecoder_toDown_d_payload_opcode = vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode;
  assign vexiis_0_iBus_noDecoder_toDown_d_payload_param = vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_param;
  assign vexiis_0_iBus_noDecoder_toDown_d_payload_denied = vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_denied;
  assign vexiis_0_iBus_noDecoder_toDown_d_payload_data = vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_data;
  assign vexiis_0_iBus_noDecoder_toDown_d_payload_corrupt = vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_corrupt;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_size = vexiis_0_iBus_noDecoder_toDown_a_payload_size;
  assign vexiis_0_iBus_noDecoder_toDown_d_payload_size = vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_size;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_address = vexiis_0_iBus_noDecoder_toDown_a_payload_address;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_valid = vexiis_0_lsuL1Bus_noDecoder_toDown_a_valid;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_a_ready = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_ready;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode = vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_opcode;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_param = vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_param;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_source = vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_source;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_mask = vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_mask;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_data = vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_data;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_corrupt = vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_corrupt;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_valid = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_valid;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_ready = vexiis_0_lsuL1Bus_noDecoder_toDown_d_ready;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_param = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_param;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_source = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_source;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_denied = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_denied;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_data = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_data;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_corrupt = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_corrupt;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_size = vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_size;
  assign vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_size = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_size;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_address = vexiis_0_lsuL1Bus_noDecoder_toDown_a_payload_address;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_valid = vexiis_0_dBus_to_ioBus_up_bus_a_valid;
  assign vexiis_0_dBus_to_ioBus_up_bus_a_ready = vexiis_0_dBus_to_ioBus_down_bus_a_ready;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode = vexiis_0_dBus_to_ioBus_up_bus_a_payload_opcode;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_payload_param = vexiis_0_dBus_to_ioBus_up_bus_a_payload_param;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_payload_address = vexiis_0_dBus_to_ioBus_up_bus_a_payload_address;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_payload_size = vexiis_0_dBus_to_ioBus_up_bus_a_payload_size;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_payload_mask = vexiis_0_dBus_to_ioBus_up_bus_a_payload_mask;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_payload_data = vexiis_0_dBus_to_ioBus_up_bus_a_payload_data;
  assign vexiis_0_dBus_to_ioBus_down_bus_a_payload_corrupt = vexiis_0_dBus_to_ioBus_up_bus_a_payload_corrupt;
  assign vexiis_0_dBus_to_ioBus_up_bus_d_valid = vexiis_0_dBus_to_ioBus_down_bus_d_valid;
  assign vexiis_0_dBus_to_ioBus_down_bus_d_ready = vexiis_0_dBus_to_ioBus_up_bus_d_ready;
  assign vexiis_0_dBus_to_ioBus_up_bus_d_payload_opcode = vexiis_0_dBus_to_ioBus_down_bus_d_payload_opcode;
  assign vexiis_0_dBus_to_ioBus_up_bus_d_payload_param = vexiis_0_dBus_to_ioBus_down_bus_d_payload_param;
  assign vexiis_0_dBus_to_ioBus_up_bus_d_payload_size = vexiis_0_dBus_to_ioBus_down_bus_d_payload_size;
  assign vexiis_0_dBus_to_ioBus_up_bus_d_payload_denied = vexiis_0_dBus_to_ioBus_down_bus_d_payload_denied;
  assign vexiis_0_dBus_to_ioBus_up_bus_d_payload_data = vexiis_0_dBus_to_ioBus_down_bus_d_payload_data;
  assign vexiis_0_dBus_to_ioBus_up_bus_d_payload_corrupt = vexiis_0_dBus_to_ioBus_down_bus_d_payload_corrupt;
  assign vexiis_0_dBus_bus_a_valid = vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_valid;
  assign vexiis_0_dBus_bus_a_payload_opcode = vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode;
  assign vexiis_0_dBus_bus_a_payload_param = vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_param;
  assign vexiis_0_dBus_bus_a_payload_address = vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_address;
  assign vexiis_0_dBus_bus_a_payload_size = vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_size;
  assign vexiis_0_dBus_bus_a_payload_mask = vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_mask;
  assign vexiis_0_dBus_bus_a_payload_data = vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_data;
  assign vexiis_0_dBus_bus_a_payload_corrupt = vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt;
  assign vexiis_0_dBus_bus_d_ready = vexiis_0_logic_core_LsuTileLinkPlugin_logic_bridge_down_d_ready;
  assign mem_toAxi4_up_bus_a_ready = mem_toAxi4_logic_bridge_io_up_a_ready;
  assign mem_toAxi4_up_bus_d_valid = mem_toAxi4_logic_bridge_io_up_d_valid;
  assign mem_toAxi4_up_bus_d_payload_opcode = mem_toAxi4_logic_bridge_io_up_d_payload_opcode;
  assign mem_toAxi4_up_bus_d_payload_param = mem_toAxi4_logic_bridge_io_up_d_payload_param;
  assign mem_toAxi4_up_bus_d_payload_source = mem_toAxi4_logic_bridge_io_up_d_payload_source;
  assign mem_toAxi4_up_bus_d_payload_size = mem_toAxi4_logic_bridge_io_up_d_payload_size;
  assign mem_toAxi4_up_bus_d_payload_denied = mem_toAxi4_logic_bridge_io_up_d_payload_denied;
  assign mem_toAxi4_up_bus_d_payload_data = mem_toAxi4_logic_bridge_io_up_d_payload_data;
  assign mem_toAxi4_up_bus_d_payload_corrupt = mem_toAxi4_logic_bridge_io_up_d_payload_corrupt;
  assign mem_toAxi4_down_ar_valid = mem_toAxi4_logic_bridge_io_down_ar_valid;
  assign mem_toAxi4_down_ar_payload_addr = mem_toAxi4_logic_bridge_io_down_ar_payload_addr;
  assign mem_toAxi4_down_ar_payload_id = mem_toAxi4_logic_bridge_io_down_ar_payload_id;
  assign mem_toAxi4_down_ar_payload_len = mem_toAxi4_logic_bridge_io_down_ar_payload_len;
  assign mem_toAxi4_down_ar_payload_size = mem_toAxi4_logic_bridge_io_down_ar_payload_size;
  assign mem_toAxi4_down_ar_payload_burst = mem_toAxi4_logic_bridge_io_down_ar_payload_burst;
  assign mem_toAxi4_down_aw_valid = mem_toAxi4_logic_bridge_io_down_aw_valid;
  assign mem_toAxi4_down_aw_payload_addr = mem_toAxi4_logic_bridge_io_down_aw_payload_addr;
  assign mem_toAxi4_down_aw_payload_id = mem_toAxi4_logic_bridge_io_down_aw_payload_id;
  assign mem_toAxi4_down_aw_payload_len = mem_toAxi4_logic_bridge_io_down_aw_payload_len;
  assign mem_toAxi4_down_aw_payload_size = mem_toAxi4_logic_bridge_io_down_aw_payload_size;
  assign mem_toAxi4_down_aw_payload_burst = mem_toAxi4_logic_bridge_io_down_aw_payload_burst;
  assign mem_toAxi4_down_aw_payload_allStrb = mem_toAxi4_logic_bridge_io_down_aw_payload_allStrb;
  assign mem_toAxi4_down_w_valid = mem_toAxi4_logic_bridge_io_down_w_valid;
  assign mem_toAxi4_down_w_payload_data = mem_toAxi4_logic_bridge_io_down_w_payload_data;
  assign mem_toAxi4_down_w_payload_strb = mem_toAxi4_logic_bridge_io_down_w_payload_strb;
  assign mem_toAxi4_down_w_payload_last = mem_toAxi4_logic_bridge_io_down_w_payload_last;
  assign mem_toAxi4_down_r_ready = mem_toAxi4_logic_bridge_io_down_r_ready;
  assign mem_toAxi4_down_b_ready = mem_toAxi4_logic_bridge_io_down_b_ready;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_a_valid = vexiis_0_iBus_to_splited_mBus_up_bus_a_valid;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_a_ready = vexiis_0_iBus_to_splited_mBus_down_bus_a_ready;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_opcode = vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_opcode;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_param = vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_param;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_address = vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_address;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_a_payload_size = vexiis_0_iBus_to_splited_mBus_up_bus_a_payload_size;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_d_valid = vexiis_0_iBus_to_splited_mBus_down_bus_d_valid;
  assign vexiis_0_iBus_to_splited_mBus_down_bus_d_ready = vexiis_0_iBus_to_splited_mBus_up_bus_d_ready;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_opcode = vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_opcode;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_param = vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_param;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_size = vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_size;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_denied = vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_denied;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_data = vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_data;
  assign vexiis_0_iBus_to_splited_mBus_up_bus_d_payload_corrupt = vexiis_0_iBus_to_splited_mBus_down_bus_d_payload_corrupt;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_valid = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_valid;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_ready = vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_ready;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_opcode = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_opcode;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_param = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_param;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_source = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_source;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_address = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_address;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_size = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_size;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_mask = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_mask;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_data = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_data;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_a_payload_corrupt = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_a_payload_corrupt;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_valid = vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_valid;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_ready = vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_ready;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_opcode = vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_opcode;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_param = vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_param;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_source = vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_source;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_size = vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_size;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_denied = vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_denied;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_data = vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_data;
  assign vexiis_0_lsuL1Bus_to_splited_mBus_up_bus_d_payload_corrupt = vexiis_0_lsuL1Bus_to_splited_mBus_down_bus_d_payload_corrupt;
  assign peripheral_clint_node_bus_a_valid = peripheral_bus_to_peripheral_clint_node_down_bus_a_valid;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_ready = peripheral_clint_node_bus_a_ready;
  assign peripheral_clint_node_bus_a_payload_opcode = peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode;
  assign peripheral_clint_node_bus_a_payload_param = peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_param;
  assign peripheral_clint_node_bus_a_payload_source = peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_source;
  assign peripheral_clint_node_bus_a_payload_address = peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_address;
  assign peripheral_clint_node_bus_a_payload_size = peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_size;
  assign peripheral_clint_node_bus_a_payload_mask = peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_mask;
  assign peripheral_clint_node_bus_a_payload_data = peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_data;
  assign peripheral_clint_node_bus_a_payload_corrupt = peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_corrupt;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_d_valid = peripheral_clint_node_bus_d_valid;
  assign peripheral_clint_node_bus_d_ready = peripheral_bus_to_peripheral_clint_node_down_bus_d_ready;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode = peripheral_clint_node_bus_d_payload_opcode;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_param = peripheral_clint_node_bus_d_payload_param;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_source = peripheral_clint_node_bus_d_payload_source;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_size = peripheral_clint_node_bus_d_payload_size;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_denied = peripheral_clint_node_bus_d_payload_denied;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_data = peripheral_clint_node_bus_d_payload_data;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_corrupt = peripheral_clint_node_bus_d_payload_corrupt;
  assign peripheral_plic_node_bus_a_valid = peripheral_bus_to_peripheral_plic_node_down_bus_a_valid;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_ready = peripheral_plic_node_bus_a_ready;
  assign peripheral_plic_node_bus_a_payload_opcode = peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode;
  assign peripheral_plic_node_bus_a_payload_param = peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_param;
  assign peripheral_plic_node_bus_a_payload_source = peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_source;
  assign peripheral_plic_node_bus_a_payload_address = peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_address;
  assign peripheral_plic_node_bus_a_payload_size = peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_size;
  assign peripheral_plic_node_bus_a_payload_mask = peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_mask;
  assign peripheral_plic_node_bus_a_payload_data = peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_data;
  assign peripheral_plic_node_bus_a_payload_corrupt = peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_corrupt;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_d_valid = peripheral_plic_node_bus_d_valid;
  assign peripheral_plic_node_bus_d_ready = peripheral_bus_to_peripheral_plic_node_down_bus_d_ready;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode = peripheral_plic_node_bus_d_payload_opcode;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_param = peripheral_plic_node_bus_d_payload_param;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_source = peripheral_plic_node_bus_d_payload_source;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_size = peripheral_plic_node_bus_d_payload_size;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_denied = peripheral_plic_node_bus_d_payload_denied;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_data = peripheral_plic_node_bus_d_payload_data;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_corrupt = peripheral_plic_node_bus_d_payload_corrupt;
  assign peripheral_toAxiLite4_up_bus_a_valid = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_valid;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_ready = peripheral_toAxiLite4_up_bus_a_ready;
  assign peripheral_toAxiLite4_up_bus_a_payload_opcode = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode;
  assign peripheral_toAxiLite4_up_bus_a_payload_param = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_param;
  assign peripheral_toAxiLite4_up_bus_a_payload_source = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_source;
  assign peripheral_toAxiLite4_up_bus_a_payload_address = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_address;
  assign peripheral_toAxiLite4_up_bus_a_payload_size = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_size;
  assign peripheral_toAxiLite4_up_bus_a_payload_mask = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_mask;
  assign peripheral_toAxiLite4_up_bus_a_payload_data = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_data;
  assign peripheral_toAxiLite4_up_bus_a_payload_corrupt = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_corrupt;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_valid = peripheral_toAxiLite4_up_bus_d_valid;
  assign peripheral_toAxiLite4_up_bus_d_ready = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_ready;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode = peripheral_toAxiLite4_up_bus_d_payload_opcode;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_param = peripheral_toAxiLite4_up_bus_d_payload_param;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_source = peripheral_toAxiLite4_up_bus_d_payload_source;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_size = peripheral_toAxiLite4_up_bus_d_payload_size;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_denied = peripheral_toAxiLite4_up_bus_d_payload_denied;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_data = peripheral_toAxiLite4_up_bus_d_payload_data;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_corrupt = peripheral_toAxiLite4_up_bus_d_payload_corrupt;
  assign ioBus_to_peripheral_bus_up_bus_a_valid = ioBus_noDecoder_toDown_a_valid;
  assign ioBus_noDecoder_toDown_a_ready = ioBus_to_peripheral_bus_up_bus_a_ready;
  assign ioBus_to_peripheral_bus_up_bus_a_payload_opcode = ioBus_noDecoder_toDown_a_payload_opcode;
  assign ioBus_to_peripheral_bus_up_bus_a_payload_param = ioBus_noDecoder_toDown_a_payload_param;
  assign ioBus_to_peripheral_bus_up_bus_a_payload_mask = ioBus_noDecoder_toDown_a_payload_mask;
  assign ioBus_to_peripheral_bus_up_bus_a_payload_data = ioBus_noDecoder_toDown_a_payload_data;
  assign ioBus_to_peripheral_bus_up_bus_a_payload_corrupt = ioBus_noDecoder_toDown_a_payload_corrupt;
  assign ioBus_noDecoder_toDown_d_valid = ioBus_to_peripheral_bus_up_bus_d_valid;
  assign ioBus_to_peripheral_bus_up_bus_d_ready = ioBus_noDecoder_toDown_d_ready;
  assign ioBus_noDecoder_toDown_d_payload_opcode = ioBus_to_peripheral_bus_up_bus_d_payload_opcode;
  assign ioBus_noDecoder_toDown_d_payload_param = ioBus_to_peripheral_bus_up_bus_d_payload_param;
  assign ioBus_noDecoder_toDown_d_payload_denied = ioBus_to_peripheral_bus_up_bus_d_payload_denied;
  assign ioBus_noDecoder_toDown_d_payload_data = ioBus_to_peripheral_bus_up_bus_d_payload_data;
  assign ioBus_noDecoder_toDown_d_payload_corrupt = ioBus_to_peripheral_bus_up_bus_d_payload_corrupt;
  assign ioBus_to_peripheral_bus_up_bus_a_payload_size = ioBus_noDecoder_toDown_a_payload_size;
  assign ioBus_noDecoder_toDown_d_payload_size = ioBus_to_peripheral_bus_up_bus_d_payload_size;
  assign ioBus_to_peripheral_bus_up_bus_a_payload_address = ioBus_noDecoder_toDown_a_payload_address;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_valid = splited_mBus_decoder_core_io_downs_0_a_valid;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_opcode = splited_mBus_decoder_core_io_downs_0_a_payload_opcode;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_param = splited_mBus_decoder_core_io_downs_0_a_payload_param;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_source = splited_mBus_decoder_core_io_downs_0_a_payload_source;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_address = splited_mBus_decoder_core_io_downs_0_a_payload_address;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_size = splited_mBus_decoder_core_io_downs_0_a_payload_size;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_mask = splited_mBus_decoder_core_io_downs_0_a_payload_mask;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_data = splited_mBus_decoder_core_io_downs_0_a_payload_data;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_payload_corrupt = splited_mBus_decoder_core_io_downs_0_a_payload_corrupt;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_d_ready = splited_mBus_decoder_core_io_downs_0_d_ready;
  assign splited_mBus_to_peripheral_bus_up_bus_a_valid = splited_mBus_decoder_core_io_downs_1_a_valid;
  assign splited_mBus_to_peripheral_bus_up_bus_a_payload_opcode = splited_mBus_decoder_core_io_downs_1_a_payload_opcode;
  assign splited_mBus_to_peripheral_bus_up_bus_a_payload_param = splited_mBus_decoder_core_io_downs_1_a_payload_param;
  assign splited_mBus_to_peripheral_bus_up_bus_a_payload_source = splited_mBus_decoder_core_io_downs_1_a_payload_source;
  assign splited_mBus_to_peripheral_bus_up_bus_a_payload_address = splited_mBus_decoder_core_io_downs_1_a_payload_address;
  assign splited_mBus_to_peripheral_bus_up_bus_a_payload_size = splited_mBus_decoder_core_io_downs_1_a_payload_size;
  assign splited_mBus_to_peripheral_bus_up_bus_a_payload_mask = splited_mBus_decoder_core_io_downs_1_a_payload_mask;
  assign splited_mBus_to_peripheral_bus_up_bus_a_payload_data = splited_mBus_decoder_core_io_downs_1_a_payload_data;
  assign splited_mBus_to_peripheral_bus_up_bus_a_payload_corrupt = splited_mBus_decoder_core_io_downs_1_a_payload_corrupt;
  assign splited_mBus_to_peripheral_bus_up_bus_d_ready = splited_mBus_decoder_core_io_downs_1_d_ready;
  assign splited_mBus_bus_a_ready = splited_mBus_decoder_core_io_up_a_ready;
  assign splited_mBus_bus_d_valid = splited_mBus_decoder_core_io_up_d_valid;
  assign splited_mBus_bus_d_payload_opcode = splited_mBus_decoder_core_io_up_d_payload_opcode;
  assign splited_mBus_bus_d_payload_param = splited_mBus_decoder_core_io_up_d_payload_param;
  assign splited_mBus_bus_d_payload_source = splited_mBus_decoder_core_io_up_d_payload_source;
  assign splited_mBus_bus_d_payload_size = splited_mBus_decoder_core_io_up_d_payload_size;
  assign splited_mBus_bus_d_payload_denied = splited_mBus_decoder_core_io_up_d_payload_denied;
  assign splited_mBus_bus_d_payload_data = splited_mBus_decoder_core_io_up_d_payload_data;
  assign splited_mBus_bus_d_payload_corrupt = splited_mBus_decoder_core_io_up_d_payload_corrupt;
  assign mBusAxi_ar_valid = mem_toAxi4_down_ar_valid;
  assign mem_toAxi4_down_ar_ready = mBusAxi_ar_ready;
  assign mBusAxi_ar_payload_addr = mem_toAxi4_down_ar_payload_addr;
  assign mBusAxi_ar_payload_id = {6'd0, mem_toAxi4_down_ar_payload_id};
  assign mBusAxi_ar_payload_len = mem_toAxi4_down_ar_payload_len;
  assign mBusAxi_ar_payload_size = mem_toAxi4_down_ar_payload_size;
  assign mBusAxi_ar_payload_burst = mem_toAxi4_down_ar_payload_burst;
  assign mBusAxi_aw_valid = mem_toAxi4_down_aw_valid;
  assign mem_toAxi4_down_aw_ready = mBusAxi_aw_ready;
  assign mBusAxi_aw_payload_addr = mem_toAxi4_down_aw_payload_addr;
  assign mBusAxi_aw_payload_id = {6'd0, mem_toAxi4_down_aw_payload_id};
  assign mBusAxi_aw_payload_len = mem_toAxi4_down_aw_payload_len;
  assign mBusAxi_aw_payload_size = mem_toAxi4_down_aw_payload_size;
  assign mBusAxi_aw_payload_burst = mem_toAxi4_down_aw_payload_burst;
  assign mBusAxi_aw_payload_allStrb = mem_toAxi4_down_aw_payload_allStrb;
  assign mBusAxi_w_valid = mem_toAxi4_down_w_valid;
  assign mem_toAxi4_down_w_ready = mBusAxi_w_ready;
  assign mBusAxi_w_payload_data = mem_toAxi4_down_w_payload_data;
  assign mBusAxi_w_payload_strb = mem_toAxi4_down_w_payload_strb;
  assign mBusAxi_w_payload_last = mem_toAxi4_down_w_payload_last;
  assign mem_toAxi4_down_r_valid = mBusAxi_r_valid;
  assign mBusAxi_r_ready = mem_toAxi4_down_r_ready;
  assign mem_toAxi4_down_r_payload_data = mBusAxi_r_payload_data;
  assign mem_toAxi4_down_r_payload_last = mBusAxi_r_payload_last;
  assign mem_toAxi4_down_r_payload_id = mBusAxi_r_payload_id[1:0];
  assign mem_toAxi4_down_r_payload_resp = mBusAxi_r_payload_resp;
  assign mem_toAxi4_down_b_valid = mBusAxi_b_valid;
  assign mBusAxi_b_ready = mem_toAxi4_down_b_ready;
  assign mem_toAxi4_down_b_payload_id = mBusAxi_b_payload_id[1:0];
  assign mem_toAxi4_down_b_payload_resp = mBusAxi_b_payload_resp;
  assign mBusAxi_aw_ready = mBusAxi_aw_rValidN;
  assign mBusAxi_aw_s2mPipe_valid = (mBusAxi_aw_valid || (! mBusAxi_aw_rValidN));
  assign mBusAxi_aw_s2mPipe_payload_addr = (mBusAxi_aw_rValidN ? mBusAxi_aw_payload_addr : mBusAxi_aw_rData_addr);
  assign mBusAxi_aw_s2mPipe_payload_id = (mBusAxi_aw_rValidN ? mBusAxi_aw_payload_id : mBusAxi_aw_rData_id);
  assign mBusAxi_aw_s2mPipe_payload_len = (mBusAxi_aw_rValidN ? mBusAxi_aw_payload_len : mBusAxi_aw_rData_len);
  assign mBusAxi_aw_s2mPipe_payload_size = (mBusAxi_aw_rValidN ? mBusAxi_aw_payload_size : mBusAxi_aw_rData_size);
  assign mBusAxi_aw_s2mPipe_payload_burst = (mBusAxi_aw_rValidN ? mBusAxi_aw_payload_burst : mBusAxi_aw_rData_burst);
  assign mBusAxi_aw_s2mPipe_payload_allStrb = (mBusAxi_aw_rValidN ? mBusAxi_aw_payload_allStrb : mBusAxi_aw_rData_allStrb);
  always @(*) begin
    mBusAxi_aw_s2mPipe_ready = mBusAxi_aw_s2mPipe_m2sPipe_ready;
    if(when_Stream_l399_4) begin
      mBusAxi_aw_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l399_4 = (! mBusAxi_aw_s2mPipe_m2sPipe_valid);
  assign mBusAxi_aw_s2mPipe_m2sPipe_valid = mBusAxi_aw_s2mPipe_rValid;
  assign mBusAxi_aw_s2mPipe_m2sPipe_payload_addr = mBusAxi_aw_s2mPipe_rData_addr;
  assign mBusAxi_aw_s2mPipe_m2sPipe_payload_id = mBusAxi_aw_s2mPipe_rData_id;
  assign mBusAxi_aw_s2mPipe_m2sPipe_payload_len = mBusAxi_aw_s2mPipe_rData_len;
  assign mBusAxi_aw_s2mPipe_m2sPipe_payload_size = mBusAxi_aw_s2mPipe_rData_size;
  assign mBusAxi_aw_s2mPipe_m2sPipe_payload_burst = mBusAxi_aw_s2mPipe_rData_burst;
  assign mBusAxi_aw_s2mPipe_m2sPipe_payload_allStrb = mBusAxi_aw_s2mPipe_rData_allStrb;
  assign mBus_awvalid = mBusAxi_aw_s2mPipe_m2sPipe_valid;
  assign mBusAxi_aw_s2mPipe_m2sPipe_ready = mBus_awready;
  assign mBus_awaddr = mBusAxi_aw_s2mPipe_m2sPipe_payload_addr;
  assign mBus_awid = mBusAxi_aw_s2mPipe_m2sPipe_payload_id;
  assign mBus_awlen = mBusAxi_aw_s2mPipe_m2sPipe_payload_len;
  assign mBus_awsize = mBusAxi_aw_s2mPipe_m2sPipe_payload_size;
  assign mBus_awburst = mBusAxi_aw_s2mPipe_m2sPipe_payload_burst;
  assign mBus_awallStrb = mBusAxi_aw_s2mPipe_m2sPipe_payload_allStrb;
  assign mBusAxi_w_ready = mBusAxi_w_rValidN;
  assign mBusAxi_w_s2mPipe_valid = (mBusAxi_w_valid || (! mBusAxi_w_rValidN));
  assign mBusAxi_w_s2mPipe_payload_data = (mBusAxi_w_rValidN ? mBusAxi_w_payload_data : mBusAxi_w_rData_data);
  assign mBusAxi_w_s2mPipe_payload_strb = (mBusAxi_w_rValidN ? mBusAxi_w_payload_strb : mBusAxi_w_rData_strb);
  assign mBusAxi_w_s2mPipe_payload_last = (mBusAxi_w_rValidN ? mBusAxi_w_payload_last : mBusAxi_w_rData_last);
  always @(*) begin
    mBusAxi_w_s2mPipe_ready = mBusAxi_w_s2mPipe_m2sPipe_ready;
    if(when_Stream_l399_5) begin
      mBusAxi_w_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l399_5 = (! mBusAxi_w_s2mPipe_m2sPipe_valid);
  assign mBusAxi_w_s2mPipe_m2sPipe_valid = mBusAxi_w_s2mPipe_rValid;
  assign mBusAxi_w_s2mPipe_m2sPipe_payload_data = mBusAxi_w_s2mPipe_rData_data;
  assign mBusAxi_w_s2mPipe_m2sPipe_payload_strb = mBusAxi_w_s2mPipe_rData_strb;
  assign mBusAxi_w_s2mPipe_m2sPipe_payload_last = mBusAxi_w_s2mPipe_rData_last;
  assign mBus_wvalid = mBusAxi_w_s2mPipe_m2sPipe_valid;
  assign mBusAxi_w_s2mPipe_m2sPipe_ready = mBus_wready;
  assign mBus_wdata = mBusAxi_w_s2mPipe_m2sPipe_payload_data;
  assign mBus_wstrb = mBusAxi_w_s2mPipe_m2sPipe_payload_strb;
  assign mBus_wlast = mBusAxi_w_s2mPipe_m2sPipe_payload_last;
  assign mBus_bready = mBus_b_rValidN;
  assign mBus_b_s2mPipe_valid = (mBus_bvalid || (! mBus_b_rValidN));
  assign mBus_b_s2mPipe_payload_id = (mBus_b_rValidN ? mBus_bid : mBus_b_rData_id);
  assign mBus_b_s2mPipe_payload_resp = (mBus_b_rValidN ? mBus_bresp : mBus_b_rData_resp);
  always @(*) begin
    mBus_b_s2mPipe_ready = mBus_b_s2mPipe_m2sPipe_ready;
    if(when_Stream_l399_6) begin
      mBus_b_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l399_6 = (! mBus_b_s2mPipe_m2sPipe_valid);
  assign mBus_b_s2mPipe_m2sPipe_valid = mBus_b_s2mPipe_rValid;
  assign mBus_b_s2mPipe_m2sPipe_payload_id = mBus_b_s2mPipe_rData_id;
  assign mBus_b_s2mPipe_m2sPipe_payload_resp = mBus_b_s2mPipe_rData_resp;
  assign mBusAxi_b_valid = mBus_b_s2mPipe_m2sPipe_valid;
  assign mBus_b_s2mPipe_m2sPipe_ready = mBusAxi_b_ready;
  assign mBusAxi_b_payload_id = mBus_b_s2mPipe_m2sPipe_payload_id;
  assign mBusAxi_b_payload_resp = mBus_b_s2mPipe_m2sPipe_payload_resp;
  assign mBusAxi_ar_ready = mBusAxi_ar_rValidN;
  assign mBusAxi_ar_s2mPipe_valid = (mBusAxi_ar_valid || (! mBusAxi_ar_rValidN));
  assign mBusAxi_ar_s2mPipe_payload_addr = (mBusAxi_ar_rValidN ? mBusAxi_ar_payload_addr : mBusAxi_ar_rData_addr);
  assign mBusAxi_ar_s2mPipe_payload_id = (mBusAxi_ar_rValidN ? mBusAxi_ar_payload_id : mBusAxi_ar_rData_id);
  assign mBusAxi_ar_s2mPipe_payload_len = (mBusAxi_ar_rValidN ? mBusAxi_ar_payload_len : mBusAxi_ar_rData_len);
  assign mBusAxi_ar_s2mPipe_payload_size = (mBusAxi_ar_rValidN ? mBusAxi_ar_payload_size : mBusAxi_ar_rData_size);
  assign mBusAxi_ar_s2mPipe_payload_burst = (mBusAxi_ar_rValidN ? mBusAxi_ar_payload_burst : mBusAxi_ar_rData_burst);
  always @(*) begin
    mBusAxi_ar_s2mPipe_ready = mBusAxi_ar_s2mPipe_m2sPipe_ready;
    if(when_Stream_l399_7) begin
      mBusAxi_ar_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l399_7 = (! mBusAxi_ar_s2mPipe_m2sPipe_valid);
  assign mBusAxi_ar_s2mPipe_m2sPipe_valid = mBusAxi_ar_s2mPipe_rValid;
  assign mBusAxi_ar_s2mPipe_m2sPipe_payload_addr = mBusAxi_ar_s2mPipe_rData_addr;
  assign mBusAxi_ar_s2mPipe_m2sPipe_payload_id = mBusAxi_ar_s2mPipe_rData_id;
  assign mBusAxi_ar_s2mPipe_m2sPipe_payload_len = mBusAxi_ar_s2mPipe_rData_len;
  assign mBusAxi_ar_s2mPipe_m2sPipe_payload_size = mBusAxi_ar_s2mPipe_rData_size;
  assign mBusAxi_ar_s2mPipe_m2sPipe_payload_burst = mBusAxi_ar_s2mPipe_rData_burst;
  assign mBus_arvalid = mBusAxi_ar_s2mPipe_m2sPipe_valid;
  assign mBusAxi_ar_s2mPipe_m2sPipe_ready = mBus_arready;
  assign mBus_araddr = mBusAxi_ar_s2mPipe_m2sPipe_payload_addr;
  assign mBus_arid = mBusAxi_ar_s2mPipe_m2sPipe_payload_id;
  assign mBus_arlen = mBusAxi_ar_s2mPipe_m2sPipe_payload_len;
  assign mBus_arsize = mBusAxi_ar_s2mPipe_m2sPipe_payload_size;
  assign mBus_arburst = mBusAxi_ar_s2mPipe_m2sPipe_payload_burst;
  assign mBus_rready = mBus_r_rValidN;
  assign mBus_r_s2mPipe_valid = (mBus_rvalid || (! mBus_r_rValidN));
  assign mBus_r_s2mPipe_payload_data = (mBus_r_rValidN ? mBus_rdata : mBus_r_rData_data);
  assign mBus_r_s2mPipe_payload_id = (mBus_r_rValidN ? mBus_rid : mBus_r_rData_id);
  assign mBus_r_s2mPipe_payload_resp = (mBus_r_rValidN ? mBus_rresp : mBus_r_rData_resp);
  assign mBus_r_s2mPipe_payload_last = (mBus_r_rValidN ? mBus_rlast : mBus_r_rData_last);
  always @(*) begin
    mBus_r_s2mPipe_ready = mBus_r_s2mPipe_m2sPipe_ready;
    if(when_Stream_l399_8) begin
      mBus_r_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l399_8 = (! mBus_r_s2mPipe_m2sPipe_valid);
  assign mBus_r_s2mPipe_m2sPipe_valid = mBus_r_s2mPipe_rValid;
  assign mBus_r_s2mPipe_m2sPipe_payload_data = mBus_r_s2mPipe_rData_data;
  assign mBus_r_s2mPipe_m2sPipe_payload_id = mBus_r_s2mPipe_rData_id;
  assign mBus_r_s2mPipe_m2sPipe_payload_resp = mBus_r_s2mPipe_rData_resp;
  assign mBus_r_s2mPipe_m2sPipe_payload_last = mBus_r_s2mPipe_rData_last;
  assign mBusAxi_r_valid = mBus_r_s2mPipe_m2sPipe_valid;
  assign mBus_r_s2mPipe_m2sPipe_ready = mBusAxi_r_ready;
  assign mBusAxi_r_payload_data = mBus_r_s2mPipe_m2sPipe_payload_data;
  assign mBusAxi_r_payload_id = mBus_r_s2mPipe_m2sPipe_payload_id;
  assign mBusAxi_r_payload_resp = mBus_r_s2mPipe_m2sPipe_payload_resp;
  assign mBusAxi_r_payload_last = mBus_r_s2mPipe_m2sPipe_payload_last;
  assign vexiis_0_cfuBus_node_cmd_valid = vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_valid;
  assign vexiis_0_cfuBus_node_rsp_ready = vexiis_0_logic_core_CfuPlugin_logic_bus_rsp_ready;
  assign vexiis_0_cfuBus_node_cmd_payload_function_id = vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_function_id;
  assign vexiis_0_cfuBus_node_cmd_payload_inputs_0 = vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_inputs_0;
  assign vexiis_0_cfuBus_node_cmd_payload_inputs_1 = vexiis_0_logic_core_CfuPlugin_logic_bus_cmd_payload_inputs_1;
  assign vexiis_0_priv_stoptime = 1'b0;
  assign peripheral_clint_node_bus_a_ready = peripheral_clint_thread_core_io_bus_a_ready;
  assign peripheral_clint_node_bus_d_valid = peripheral_clint_thread_core_io_bus_d_valid;
  assign peripheral_clint_node_bus_d_payload_opcode = peripheral_clint_thread_core_io_bus_d_payload_opcode;
  assign peripheral_clint_node_bus_d_payload_param = peripheral_clint_thread_core_io_bus_d_payload_param;
  assign peripheral_clint_node_bus_d_payload_source = peripheral_clint_thread_core_io_bus_d_payload_source;
  assign peripheral_clint_node_bus_d_payload_size = peripheral_clint_thread_core_io_bus_d_payload_size;
  assign peripheral_clint_node_bus_d_payload_denied = peripheral_clint_thread_core_io_bus_d_payload_denied;
  assign peripheral_clint_node_bus_d_payload_data = peripheral_clint_thread_core_io_bus_d_payload_data;
  assign peripheral_clint_node_bus_d_payload_corrupt = peripheral_clint_thread_core_io_bus_d_payload_corrupt;
  assign peripheral_clint_thread_core_io_stop = (&vexiis_0_priv_stoptime_regNext);
  assign peripheral_clint_time = peripheral_clint_thread_core_io_time;
  assign peripheral_plic_node_bus_a_ready = peripheral_plic_thread_logic_io_bus_a_ready;
  assign peripheral_plic_node_bus_d_valid = peripheral_plic_thread_logic_io_bus_d_valid;
  assign peripheral_plic_node_bus_d_payload_opcode = peripheral_plic_thread_logic_io_bus_d_payload_opcode;
  assign peripheral_plic_node_bus_d_payload_param = peripheral_plic_thread_logic_io_bus_d_payload_param;
  assign peripheral_plic_node_bus_d_payload_source = peripheral_plic_thread_logic_io_bus_d_payload_source;
  assign peripheral_plic_node_bus_d_payload_size = peripheral_plic_thread_logic_io_bus_d_payload_size;
  assign peripheral_plic_node_bus_d_payload_denied = peripheral_plic_thread_logic_io_bus_d_payload_denied;
  assign peripheral_plic_node_bus_d_payload_data = peripheral_plic_thread_logic_io_bus_d_payload_data;
  assign peripheral_plic_node_bus_d_payload_corrupt = peripheral_plic_thread_logic_io_bus_d_payload_corrupt;
  always @(*) begin
    peripheral_plic_thread_logic_io_sources[0] = peripheral_externalInterrupts_toPlic_1_node_flag;
    peripheral_plic_thread_logic_io_sources[1] = peripheral_externalInterrupts_toPlic_2_node_flag;
    peripheral_plic_thread_logic_io_sources[2] = peripheral_externalInterrupts_toPlic_3_node_flag;
    peripheral_plic_thread_logic_io_sources[3] = peripheral_externalInterrupts_toPlic_4_node_flag;
    peripheral_plic_thread_logic_io_sources[4] = peripheral_externalInterrupts_toPlic_5_node_flag;
    peripheral_plic_thread_logic_io_sources[5] = peripheral_externalInterrupts_toPlic_6_node_flag;
    peripheral_plic_thread_logic_io_sources[6] = peripheral_externalInterrupts_toPlic_7_node_flag;
    peripheral_plic_thread_logic_io_sources[7] = peripheral_externalInterrupts_toPlic_8_node_flag;
    peripheral_plic_thread_logic_io_sources[8] = peripheral_externalInterrupts_toPlic_9_node_flag;
    peripheral_plic_thread_logic_io_sources[9] = peripheral_externalInterrupts_toPlic_10_node_flag;
    peripheral_plic_thread_logic_io_sources[10] = peripheral_externalInterrupts_toPlic_11_node_flag;
    peripheral_plic_thread_logic_io_sources[11] = peripheral_externalInterrupts_toPlic_12_node_flag;
    peripheral_plic_thread_logic_io_sources[12] = peripheral_externalInterrupts_toPlic_13_node_flag;
    peripheral_plic_thread_logic_io_sources[13] = peripheral_externalInterrupts_toPlic_14_node_flag;
    peripheral_plic_thread_logic_io_sources[14] = peripheral_externalInterrupts_toPlic_15_node_flag;
    peripheral_plic_thread_logic_io_sources[15] = peripheral_externalInterrupts_toPlic_16_node_flag;
    peripheral_plic_thread_logic_io_sources[16] = peripheral_externalInterrupts_toPlic_17_node_flag;
    peripheral_plic_thread_logic_io_sources[17] = peripheral_externalInterrupts_toPlic_18_node_flag;
    peripheral_plic_thread_logic_io_sources[18] = peripheral_externalInterrupts_toPlic_19_node_flag;
    peripheral_plic_thread_logic_io_sources[19] = peripheral_externalInterrupts_toPlic_20_node_flag;
    peripheral_plic_thread_logic_io_sources[20] = peripheral_externalInterrupts_toPlic_21_node_flag;
    peripheral_plic_thread_logic_io_sources[21] = peripheral_externalInterrupts_toPlic_22_node_flag;
    peripheral_plic_thread_logic_io_sources[22] = peripheral_externalInterrupts_toPlic_23_node_flag;
    peripheral_plic_thread_logic_io_sources[23] = peripheral_externalInterrupts_toPlic_24_node_flag;
    peripheral_plic_thread_logic_io_sources[24] = peripheral_externalInterrupts_toPlic_25_node_flag;
    peripheral_plic_thread_logic_io_sources[25] = peripheral_externalInterrupts_toPlic_26_node_flag;
    peripheral_plic_thread_logic_io_sources[26] = peripheral_externalInterrupts_toPlic_27_node_flag;
    peripheral_plic_thread_logic_io_sources[27] = peripheral_externalInterrupts_toPlic_28_node_flag;
    peripheral_plic_thread_logic_io_sources[28] = peripheral_externalInterrupts_toPlic_29_node_flag;
    peripheral_plic_thread_logic_io_sources[29] = peripheral_externalInterrupts_toPlic_30_node_flag;
    peripheral_plic_thread_logic_io_sources[30] = peripheral_externalInterrupts_toPlic_31_node_flag;
  end

  assign peripheral_plic_to_vexiis_0_priv_mei_flag = peripheral_plic_thread_logic_io_targets[0];
  assign peripheral_plic_to_vexiis_0_priv_sei_flag = peripheral_plic_thread_logic_io_targets[1];
  assign peripheral_toAxiLite4_up_bus_a_ready = peripheral_toAxiLite4_logic_bridge_io_up_a_ready;
  assign peripheral_toAxiLite4_up_bus_d_valid = peripheral_toAxiLite4_logic_bridge_io_up_d_valid;
  assign peripheral_toAxiLite4_up_bus_d_payload_opcode = peripheral_toAxiLite4_logic_bridge_io_up_d_payload_opcode;
  assign peripheral_toAxiLite4_up_bus_d_payload_param = peripheral_toAxiLite4_logic_bridge_io_up_d_payload_param;
  assign peripheral_toAxiLite4_up_bus_d_payload_source = peripheral_toAxiLite4_logic_bridge_io_up_d_payload_source;
  assign peripheral_toAxiLite4_up_bus_d_payload_size = peripheral_toAxiLite4_logic_bridge_io_up_d_payload_size;
  assign peripheral_toAxiLite4_up_bus_d_payload_denied = peripheral_toAxiLite4_logic_bridge_io_up_d_payload_denied;
  assign peripheral_toAxiLite4_up_bus_d_payload_data = peripheral_toAxiLite4_logic_bridge_io_up_d_payload_data;
  assign peripheral_toAxiLite4_up_bus_d_payload_corrupt = peripheral_toAxiLite4_logic_bridge_io_up_d_payload_corrupt;
  assign peripheral_toAxiLite4_down_aw_valid = peripheral_toAxiLite4_logic_bridge_io_down_aw_valid;
  assign peripheral_toAxiLite4_down_aw_payload_addr = peripheral_toAxiLite4_logic_bridge_io_down_aw_payload_addr;
  assign peripheral_toAxiLite4_down_aw_payload_prot = peripheral_toAxiLite4_logic_bridge_io_down_aw_payload_prot;
  assign peripheral_toAxiLite4_down_w_valid = peripheral_toAxiLite4_logic_bridge_io_down_w_valid;
  assign peripheral_toAxiLite4_down_w_payload_data = peripheral_toAxiLite4_logic_bridge_io_down_w_payload_data;
  assign peripheral_toAxiLite4_down_w_payload_strb = peripheral_toAxiLite4_logic_bridge_io_down_w_payload_strb;
  assign peripheral_toAxiLite4_down_b_ready = peripheral_toAxiLite4_logic_bridge_io_down_b_ready;
  assign peripheral_toAxiLite4_down_ar_valid = peripheral_toAxiLite4_logic_bridge_io_down_ar_valid;
  assign peripheral_toAxiLite4_down_ar_payload_addr = peripheral_toAxiLite4_logic_bridge_io_down_ar_payload_addr;
  assign peripheral_toAxiLite4_down_ar_payload_prot = peripheral_toAxiLite4_logic_bridge_io_down_ar_payload_prot;
  assign peripheral_toAxiLite4_down_r_ready = peripheral_toAxiLite4_logic_bridge_io_down_r_ready;
  assign ioBus_to_peripheral_bus_down_bus_a_valid = ioBus_to_peripheral_bus_up_bus_a_valid;
  assign ioBus_to_peripheral_bus_up_bus_a_ready = ioBus_to_peripheral_bus_down_bus_a_ready;
  assign ioBus_to_peripheral_bus_down_bus_a_payload_opcode = ioBus_to_peripheral_bus_up_bus_a_payload_opcode;
  assign ioBus_to_peripheral_bus_down_bus_a_payload_param = ioBus_to_peripheral_bus_up_bus_a_payload_param;
  assign ioBus_to_peripheral_bus_down_bus_a_payload_address = ioBus_to_peripheral_bus_up_bus_a_payload_address;
  assign ioBus_to_peripheral_bus_down_bus_a_payload_size = ioBus_to_peripheral_bus_up_bus_a_payload_size;
  assign ioBus_to_peripheral_bus_down_bus_a_payload_mask = ioBus_to_peripheral_bus_up_bus_a_payload_mask;
  assign ioBus_to_peripheral_bus_down_bus_a_payload_data = ioBus_to_peripheral_bus_up_bus_a_payload_data;
  assign ioBus_to_peripheral_bus_down_bus_a_payload_corrupt = ioBus_to_peripheral_bus_up_bus_a_payload_corrupt;
  assign ioBus_to_peripheral_bus_up_bus_d_valid = ioBus_to_peripheral_bus_down_bus_d_valid;
  assign ioBus_to_peripheral_bus_down_bus_d_ready = ioBus_to_peripheral_bus_up_bus_d_ready;
  assign ioBus_to_peripheral_bus_up_bus_d_payload_opcode = ioBus_to_peripheral_bus_down_bus_d_payload_opcode;
  assign ioBus_to_peripheral_bus_up_bus_d_payload_param = ioBus_to_peripheral_bus_down_bus_d_payload_param;
  assign ioBus_to_peripheral_bus_up_bus_d_payload_size = ioBus_to_peripheral_bus_down_bus_d_payload_size;
  assign ioBus_to_peripheral_bus_up_bus_d_payload_denied = ioBus_to_peripheral_bus_down_bus_d_payload_denied;
  assign ioBus_to_peripheral_bus_up_bus_d_payload_data = ioBus_to_peripheral_bus_down_bus_d_payload_data;
  assign ioBus_to_peripheral_bus_up_bus_d_payload_corrupt = ioBus_to_peripheral_bus_down_bus_d_payload_corrupt;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_a_ready = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_a_ready;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_d_valid = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_valid;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_opcode = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_opcode;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_param = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_param;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_source = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_source;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_size = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_size;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_denied = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_denied;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_data = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_data;
  assign splited_mBus_to_mem_toAxi4_up_up_bus_d_payload_corrupt = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_up_d_payload_corrupt;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_valid = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_valid;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_opcode = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_opcode;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_param = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_param;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_source = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_source;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_address = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_address;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_size = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_size;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_mask = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_mask;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_data = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_data;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_a_payload_corrupt = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_a_payload_corrupt;
  assign splited_mBus_to_mem_toAxi4_up_down_bus_d_ready = splited_mBus_to_mem_toAxi4_up_widthAdapter_io_down_d_ready;
  assign splited_mBus_to_peripheral_bus_up_bus_a_ready = splited_mBus_to_peripheral_bus_widthAdapter_io_up_a_ready;
  assign splited_mBus_to_peripheral_bus_up_bus_d_valid = splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_valid;
  assign splited_mBus_to_peripheral_bus_up_bus_d_payload_opcode = splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_opcode;
  assign splited_mBus_to_peripheral_bus_up_bus_d_payload_param = splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_param;
  assign splited_mBus_to_peripheral_bus_up_bus_d_payload_source = splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_source;
  assign splited_mBus_to_peripheral_bus_up_bus_d_payload_size = splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_size;
  assign splited_mBus_to_peripheral_bus_up_bus_d_payload_denied = splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_denied;
  assign splited_mBus_to_peripheral_bus_up_bus_d_payload_data = splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_data;
  assign splited_mBus_to_peripheral_bus_up_bus_d_payload_corrupt = splited_mBus_to_peripheral_bus_widthAdapter_io_up_d_payload_corrupt;
  assign splited_mBus_to_peripheral_bus_down_bus_a_valid = splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_valid;
  assign splited_mBus_to_peripheral_bus_down_bus_a_payload_opcode = splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_opcode;
  assign splited_mBus_to_peripheral_bus_down_bus_a_payload_param = splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_param;
  assign splited_mBus_to_peripheral_bus_down_bus_a_payload_source = splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_source;
  assign splited_mBus_to_peripheral_bus_down_bus_a_payload_address = splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_address;
  assign splited_mBus_to_peripheral_bus_down_bus_a_payload_size = splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_size;
  assign splited_mBus_to_peripheral_bus_down_bus_a_payload_mask = splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_mask;
  assign splited_mBus_to_peripheral_bus_down_bus_a_payload_data = splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_data;
  assign splited_mBus_to_peripheral_bus_down_bus_a_payload_corrupt = splited_mBus_to_peripheral_bus_widthAdapter_io_down_a_payload_corrupt;
  assign splited_mBus_to_peripheral_bus_down_bus_d_ready = splited_mBus_to_peripheral_bus_widthAdapter_io_down_d_ready;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_valid = peripheral_bus_decoder_core_io_downs_0_a_valid;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode = peripheral_bus_decoder_core_io_downs_0_a_payload_opcode;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_param = peripheral_bus_decoder_core_io_downs_0_a_payload_param;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_source = peripheral_bus_decoder_core_io_downs_0_a_payload_source;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_address = peripheral_bus_decoder_core_io_downs_0_a_payload_address;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_size = peripheral_bus_decoder_core_io_downs_0_a_payload_size;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_mask = peripheral_bus_decoder_core_io_downs_0_a_payload_mask;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_data = peripheral_bus_decoder_core_io_downs_0_a_payload_data;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_corrupt = peripheral_bus_decoder_core_io_downs_0_a_payload_corrupt;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_d_ready = peripheral_bus_decoder_core_io_downs_0_d_ready;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_valid = peripheral_bus_decoder_core_io_downs_1_a_valid;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode = peripheral_bus_decoder_core_io_downs_1_a_payload_opcode;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_param = peripheral_bus_decoder_core_io_downs_1_a_payload_param;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_source = peripheral_bus_decoder_core_io_downs_1_a_payload_source;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_address = peripheral_bus_decoder_core_io_downs_1_a_payload_address;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_size = peripheral_bus_decoder_core_io_downs_1_a_payload_size;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_mask = peripheral_bus_decoder_core_io_downs_1_a_payload_mask;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_data = peripheral_bus_decoder_core_io_downs_1_a_payload_data;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_corrupt = peripheral_bus_decoder_core_io_downs_1_a_payload_corrupt;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_d_ready = peripheral_bus_decoder_core_io_downs_1_d_ready;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_valid = peripheral_bus_decoder_core_io_downs_2_a_valid;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode = peripheral_bus_decoder_core_io_downs_2_a_payload_opcode;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_param = peripheral_bus_decoder_core_io_downs_2_a_payload_param;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_source = peripheral_bus_decoder_core_io_downs_2_a_payload_source;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_address = peripheral_bus_decoder_core_io_downs_2_a_payload_address;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_size = peripheral_bus_decoder_core_io_downs_2_a_payload_size;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_mask = peripheral_bus_decoder_core_io_downs_2_a_payload_mask;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_data = peripheral_bus_decoder_core_io_downs_2_a_payload_data;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_corrupt = peripheral_bus_decoder_core_io_downs_2_a_payload_corrupt;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_ready = peripheral_bus_decoder_core_io_downs_2_d_ready;
  assign peripheral_bus_bus_a_halfPipe_fire = (peripheral_bus_bus_a_halfPipe_valid && peripheral_bus_bus_a_halfPipe_ready);
  assign peripheral_bus_bus_a_ready = (! peripheral_bus_bus_a_rValid);
  assign peripheral_bus_bus_a_halfPipe_valid = peripheral_bus_bus_a_rValid;
  assign peripheral_bus_bus_a_halfPipe_payload_opcode = peripheral_bus_bus_a_rData_opcode;
  assign peripheral_bus_bus_a_halfPipe_payload_param = peripheral_bus_bus_a_rData_param;
  assign peripheral_bus_bus_a_halfPipe_payload_source = peripheral_bus_bus_a_rData_source;
  assign peripheral_bus_bus_a_halfPipe_payload_address = peripheral_bus_bus_a_rData_address;
  assign peripheral_bus_bus_a_halfPipe_payload_size = peripheral_bus_bus_a_rData_size;
  assign peripheral_bus_bus_a_halfPipe_payload_mask = peripheral_bus_bus_a_rData_mask;
  assign peripheral_bus_bus_a_halfPipe_payload_data = peripheral_bus_bus_a_rData_data;
  assign peripheral_bus_bus_a_halfPipe_payload_corrupt = peripheral_bus_bus_a_rData_corrupt;
  assign peripheral_bus_bus_a_halfPipe_ready = peripheral_bus_decoder_core_io_up_a_ready;
  assign io_up_d_halfPipe_fire = (io_up_d_halfPipe_valid && io_up_d_halfPipe_ready);
  assign peripheral_bus_decoder_core_io_up_d_ready = (! io_up_d_rValid);
  assign io_up_d_halfPipe_valid = io_up_d_rValid;
  assign io_up_d_halfPipe_payload_opcode = io_up_d_rData_opcode;
  assign io_up_d_halfPipe_payload_param = io_up_d_rData_param;
  assign io_up_d_halfPipe_payload_source = io_up_d_rData_source;
  assign io_up_d_halfPipe_payload_size = io_up_d_rData_size;
  assign io_up_d_halfPipe_payload_denied = io_up_d_rData_denied;
  assign io_up_d_halfPipe_payload_data = io_up_d_rData_data;
  assign io_up_d_halfPipe_payload_corrupt = io_up_d_rData_corrupt;
  assign peripheral_bus_bus_d_valid = io_up_d_halfPipe_valid;
  assign io_up_d_halfPipe_ready = peripheral_bus_bus_d_ready;
  assign peripheral_bus_bus_d_payload_opcode = io_up_d_halfPipe_payload_opcode;
  assign peripheral_bus_bus_d_payload_param = io_up_d_halfPipe_payload_param;
  assign peripheral_bus_bus_d_payload_source = io_up_d_halfPipe_payload_source;
  assign peripheral_bus_bus_d_payload_size = io_up_d_halfPipe_payload_size;
  assign peripheral_bus_bus_d_payload_denied = io_up_d_halfPipe_payload_denied;
  assign peripheral_bus_bus_d_payload_data = io_up_d_halfPipe_payload_data;
  assign peripheral_bus_bus_d_payload_corrupt = io_up_d_halfPipe_payload_corrupt;
  assign peripheral_toAxiLite4_down_aw_halfPipe_fire = (peripheral_toAxiLite4_down_aw_halfPipe_valid && peripheral_toAxiLite4_down_aw_halfPipe_ready);
  assign peripheral_toAxiLite4_down_aw_ready = (! peripheral_toAxiLite4_down_aw_rValid);
  assign peripheral_toAxiLite4_down_aw_halfPipe_valid = peripheral_toAxiLite4_down_aw_rValid;
  assign peripheral_toAxiLite4_down_aw_halfPipe_payload_addr = peripheral_toAxiLite4_down_aw_rData_addr;
  assign peripheral_toAxiLite4_down_aw_halfPipe_payload_prot = peripheral_toAxiLite4_down_aw_rData_prot;
  assign pBus_awvalid = peripheral_toAxiLite4_down_aw_halfPipe_valid;
  assign peripheral_toAxiLite4_down_aw_halfPipe_ready = pBus_awready;
  assign pBus_awaddr = peripheral_toAxiLite4_down_aw_halfPipe_payload_addr;
  assign pBus_awprot = peripheral_toAxiLite4_down_aw_halfPipe_payload_prot;
  assign peripheral_toAxiLite4_down_w_halfPipe_fire = (peripheral_toAxiLite4_down_w_halfPipe_valid && peripheral_toAxiLite4_down_w_halfPipe_ready);
  assign peripheral_toAxiLite4_down_w_ready = (! peripheral_toAxiLite4_down_w_rValid);
  assign peripheral_toAxiLite4_down_w_halfPipe_valid = peripheral_toAxiLite4_down_w_rValid;
  assign peripheral_toAxiLite4_down_w_halfPipe_payload_data = peripheral_toAxiLite4_down_w_rData_data;
  assign peripheral_toAxiLite4_down_w_halfPipe_payload_strb = peripheral_toAxiLite4_down_w_rData_strb;
  assign pBus_wvalid = peripheral_toAxiLite4_down_w_halfPipe_valid;
  assign peripheral_toAxiLite4_down_w_halfPipe_ready = pBus_wready;
  assign pBus_wdata = peripheral_toAxiLite4_down_w_halfPipe_payload_data;
  assign pBus_wstrb = peripheral_toAxiLite4_down_w_halfPipe_payload_strb;
  assign pBus_b_halfPipe_fire = (pBus_b_halfPipe_valid && pBus_b_halfPipe_ready);
  assign pBus_bready = (! pBus_b_rValid);
  assign pBus_b_halfPipe_valid = pBus_b_rValid;
  assign pBus_b_halfPipe_payload_resp = pBus_b_rData_resp;
  assign peripheral_toAxiLite4_down_b_valid = pBus_b_halfPipe_valid;
  assign pBus_b_halfPipe_ready = peripheral_toAxiLite4_down_b_ready;
  assign peripheral_toAxiLite4_down_b_payload_resp = pBus_b_halfPipe_payload_resp;
  assign peripheral_toAxiLite4_down_ar_halfPipe_fire = (peripheral_toAxiLite4_down_ar_halfPipe_valid && peripheral_toAxiLite4_down_ar_halfPipe_ready);
  assign peripheral_toAxiLite4_down_ar_ready = (! peripheral_toAxiLite4_down_ar_rValid);
  assign peripheral_toAxiLite4_down_ar_halfPipe_valid = peripheral_toAxiLite4_down_ar_rValid;
  assign peripheral_toAxiLite4_down_ar_halfPipe_payload_addr = peripheral_toAxiLite4_down_ar_rData_addr;
  assign peripheral_toAxiLite4_down_ar_halfPipe_payload_prot = peripheral_toAxiLite4_down_ar_rData_prot;
  assign pBus_arvalid = peripheral_toAxiLite4_down_ar_halfPipe_valid;
  assign peripheral_toAxiLite4_down_ar_halfPipe_ready = pBus_arready;
  assign pBus_araddr = peripheral_toAxiLite4_down_ar_halfPipe_payload_addr;
  assign pBus_arprot = peripheral_toAxiLite4_down_ar_halfPipe_payload_prot;
  assign pBus_r_halfPipe_fire = (pBus_r_halfPipe_valid && pBus_r_halfPipe_ready);
  assign pBus_rready = (! pBus_r_rValid);
  assign pBus_r_halfPipe_valid = pBus_r_rValid;
  assign pBus_r_halfPipe_payload_data = pBus_r_rData_data;
  assign pBus_r_halfPipe_payload_resp = pBus_r_rData_resp;
  assign peripheral_toAxiLite4_down_r_valid = pBus_r_halfPipe_valid;
  assign pBus_r_halfPipe_ready = peripheral_toAxiLite4_down_r_ready;
  assign peripheral_toAxiLite4_down_r_payload_data = pBus_r_halfPipe_payload_data;
  assign peripheral_toAxiLite4_down_r_payload_resp = pBus_r_halfPipe_payload_resp;
  assign debugIn = 8'h0;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_valid = peripheral_bus_to_peripheral_clint_node_up_bus_a_valid;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_a_ready = peripheral_bus_to_peripheral_clint_node_down_bus_a_ready;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_opcode = peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_opcode;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_param = peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_param;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_source = peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_source;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_address = peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_address;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_size = peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_size;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_mask = peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_mask;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_data = peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_data;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_a_payload_corrupt = peripheral_bus_to_peripheral_clint_node_up_bus_a_payload_corrupt;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_d_valid = peripheral_bus_to_peripheral_clint_node_down_bus_d_valid;
  assign peripheral_bus_to_peripheral_clint_node_down_bus_d_ready = peripheral_bus_to_peripheral_clint_node_up_bus_d_ready;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_opcode = peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_opcode;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_param = peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_param;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_source = peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_source;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_size = peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_size;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_denied = peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_denied;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_data = peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_data;
  assign peripheral_bus_to_peripheral_clint_node_up_bus_d_payload_corrupt = peripheral_bus_to_peripheral_clint_node_down_bus_d_payload_corrupt;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_valid = peripheral_bus_to_peripheral_plic_node_up_bus_a_valid;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_a_ready = peripheral_bus_to_peripheral_plic_node_down_bus_a_ready;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_opcode = peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_opcode;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_param = peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_param;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_source = peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_source;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_address = peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_address;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_size = peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_size;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_mask = peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_mask;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_data = peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_data;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_a_payload_corrupt = peripheral_bus_to_peripheral_plic_node_up_bus_a_payload_corrupt;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_d_valid = peripheral_bus_to_peripheral_plic_node_down_bus_d_valid;
  assign peripheral_bus_to_peripheral_plic_node_down_bus_d_ready = peripheral_bus_to_peripheral_plic_node_up_bus_d_ready;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_opcode = peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_opcode;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_param = peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_param;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_source = peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_source;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_size = peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_size;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_denied = peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_denied;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_data = peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_data;
  assign peripheral_bus_to_peripheral_plic_node_up_bus_d_payload_corrupt = peripheral_bus_to_peripheral_plic_node_down_bus_d_payload_corrupt;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_valid = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_valid;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_ready = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_ready;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_opcode = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_opcode;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_param = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_param;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_source = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_source;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_address = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_address;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_size = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_size;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_mask = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_mask;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_data = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_data;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_a_payload_corrupt = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_a_payload_corrupt;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_valid = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_valid;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_ready = peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_ready;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_opcode = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_opcode;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_param = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_param;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_source = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_source;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_size = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_size;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_denied = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_denied;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_data = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_data;
  assign peripheral_bus_to_peripheral_toAxiLite4_up_up_bus_d_payload_corrupt = peripheral_bus_to_peripheral_toAxiLite4_up_down_bus_d_payload_corrupt;
  always @(posedge litex_clk) begin
    vexiis_0_priv_stoptime_regNext <= vexiis_0_priv_stoptime;
    _zz_vexiis_0_priv_rdtime <= peripheral_clint_time;
    if(vexiis_0_dBus_bus_a_ready) begin
      vexiis_0_dBus_bus_a_rData_opcode <= vexiis_0_dBus_bus_a_payload_opcode;
      vexiis_0_dBus_bus_a_rData_param <= vexiis_0_dBus_bus_a_payload_param;
      vexiis_0_dBus_bus_a_rData_address <= vexiis_0_dBus_bus_a_payload_address;
      vexiis_0_dBus_bus_a_rData_size <= vexiis_0_dBus_bus_a_payload_size;
      vexiis_0_dBus_bus_a_rData_mask <= vexiis_0_dBus_bus_a_payload_mask;
      vexiis_0_dBus_bus_a_rData_data <= vexiis_0_dBus_bus_a_payload_data;
      vexiis_0_dBus_bus_a_rData_corrupt <= vexiis_0_dBus_bus_a_payload_corrupt;
    end
    if(vexiis_0_dBus_noDecoder_toDown_d_ready) begin
      vexiis_0_dBus_noDecoder_toDown_d_rData_opcode <= vexiis_0_dBus_noDecoder_toDown_d_payload_opcode;
      vexiis_0_dBus_noDecoder_toDown_d_rData_param <= vexiis_0_dBus_noDecoder_toDown_d_payload_param;
      vexiis_0_dBus_noDecoder_toDown_d_rData_size <= vexiis_0_dBus_noDecoder_toDown_d_payload_size;
      vexiis_0_dBus_noDecoder_toDown_d_rData_denied <= vexiis_0_dBus_noDecoder_toDown_d_payload_denied;
      vexiis_0_dBus_noDecoder_toDown_d_rData_data <= vexiis_0_dBus_noDecoder_toDown_d_payload_data;
      vexiis_0_dBus_noDecoder_toDown_d_rData_corrupt <= vexiis_0_dBus_noDecoder_toDown_d_payload_corrupt;
    end
    if(vexiis_0_iBus_bus_a_ready) begin
      vexiis_0_iBus_bus_a_rData_opcode <= vexiis_0_iBus_bus_a_payload_opcode;
      vexiis_0_iBus_bus_a_rData_param <= vexiis_0_iBus_bus_a_payload_param;
      vexiis_0_iBus_bus_a_rData_address <= vexiis_0_iBus_bus_a_payload_address;
      vexiis_0_iBus_bus_a_rData_size <= vexiis_0_iBus_bus_a_payload_size;
    end
    if(vexiis_0_iBus_bus_a_halfPipe_ready) begin
      vexiis_0_iBus_bus_a_halfPipe_rData_opcode <= vexiis_0_iBus_bus_a_halfPipe_payload_opcode;
      vexiis_0_iBus_bus_a_halfPipe_rData_param <= vexiis_0_iBus_bus_a_halfPipe_payload_param;
      vexiis_0_iBus_bus_a_halfPipe_rData_address <= vexiis_0_iBus_bus_a_halfPipe_payload_address;
      vexiis_0_iBus_bus_a_halfPipe_rData_size <= vexiis_0_iBus_bus_a_halfPipe_payload_size;
    end
    if(vexiis_0_iBus_noDecoder_toDown_d_ready) begin
      vexiis_0_iBus_noDecoder_toDown_d_rData_opcode <= vexiis_0_iBus_noDecoder_toDown_d_payload_opcode;
      vexiis_0_iBus_noDecoder_toDown_d_rData_param <= vexiis_0_iBus_noDecoder_toDown_d_payload_param;
      vexiis_0_iBus_noDecoder_toDown_d_rData_size <= vexiis_0_iBus_noDecoder_toDown_d_payload_size;
      vexiis_0_iBus_noDecoder_toDown_d_rData_denied <= vexiis_0_iBus_noDecoder_toDown_d_payload_denied;
      vexiis_0_iBus_noDecoder_toDown_d_rData_data <= vexiis_0_iBus_noDecoder_toDown_d_payload_data;
      vexiis_0_iBus_noDecoder_toDown_d_rData_corrupt <= vexiis_0_iBus_noDecoder_toDown_d_payload_corrupt;
    end
    if(vexiis_0_lsuL1Bus_bus_a_ready) begin
      vexiis_0_lsuL1Bus_bus_a_rData_opcode <= vexiis_0_lsuL1Bus_bus_a_payload_opcode;
      vexiis_0_lsuL1Bus_bus_a_rData_param <= vexiis_0_lsuL1Bus_bus_a_payload_param;
      vexiis_0_lsuL1Bus_bus_a_rData_source <= vexiis_0_lsuL1Bus_bus_a_payload_source;
      vexiis_0_lsuL1Bus_bus_a_rData_address <= vexiis_0_lsuL1Bus_bus_a_payload_address;
      vexiis_0_lsuL1Bus_bus_a_rData_size <= vexiis_0_lsuL1Bus_bus_a_payload_size;
      vexiis_0_lsuL1Bus_bus_a_rData_mask <= vexiis_0_lsuL1Bus_bus_a_payload_mask;
      vexiis_0_lsuL1Bus_bus_a_rData_data <= vexiis_0_lsuL1Bus_bus_a_payload_data;
      vexiis_0_lsuL1Bus_bus_a_rData_corrupt <= vexiis_0_lsuL1Bus_bus_a_payload_corrupt;
    end
    if(vexiis_0_lsuL1Bus_bus_a_s2mPipe_ready) begin
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_opcode <= vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_opcode;
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_param <= vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_param;
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_source <= vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_source;
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_address <= vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_address;
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_size <= vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_size;
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_mask <= vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_mask;
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_data <= vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_data;
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_rData_corrupt <= vexiis_0_lsuL1Bus_bus_a_s2mPipe_payload_corrupt;
    end
    if(vexiis_0_lsuL1Bus_noDecoder_toDown_d_ready) begin
      vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_opcode <= vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_opcode;
      vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_param <= vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_param;
      vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_source <= vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_source;
      vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_size <= vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_size;
      vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_denied <= vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_denied;
      vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_data <= vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_data;
      vexiis_0_lsuL1Bus_noDecoder_toDown_d_rData_corrupt <= vexiis_0_lsuL1Bus_noDecoder_toDown_d_payload_corrupt;
    end
    if(vexiis_0_dBus_to_ioBus_down_bus_a_ready) begin
      vexiis_0_dBus_to_ioBus_down_bus_a_rData_opcode <= vexiis_0_dBus_to_ioBus_down_bus_a_payload_opcode;
      vexiis_0_dBus_to_ioBus_down_bus_a_rData_param <= vexiis_0_dBus_to_ioBus_down_bus_a_payload_param;
      vexiis_0_dBus_to_ioBus_down_bus_a_rData_address <= vexiis_0_dBus_to_ioBus_down_bus_a_payload_address;
      vexiis_0_dBus_to_ioBus_down_bus_a_rData_size <= vexiis_0_dBus_to_ioBus_down_bus_a_payload_size;
      vexiis_0_dBus_to_ioBus_down_bus_a_rData_mask <= vexiis_0_dBus_to_ioBus_down_bus_a_payload_mask;
      vexiis_0_dBus_to_ioBus_down_bus_a_rData_data <= vexiis_0_dBus_to_ioBus_down_bus_a_payload_data;
      vexiis_0_dBus_to_ioBus_down_bus_a_rData_corrupt <= vexiis_0_dBus_to_ioBus_down_bus_a_payload_corrupt;
    end
    if(mBusAxi_aw_ready) begin
      mBusAxi_aw_rData_addr <= mBusAxi_aw_payload_addr;
      mBusAxi_aw_rData_id <= mBusAxi_aw_payload_id;
      mBusAxi_aw_rData_len <= mBusAxi_aw_payload_len;
      mBusAxi_aw_rData_size <= mBusAxi_aw_payload_size;
      mBusAxi_aw_rData_burst <= mBusAxi_aw_payload_burst;
      mBusAxi_aw_rData_allStrb <= mBusAxi_aw_payload_allStrb;
    end
    if(mBusAxi_aw_s2mPipe_ready) begin
      mBusAxi_aw_s2mPipe_rData_addr <= mBusAxi_aw_s2mPipe_payload_addr;
      mBusAxi_aw_s2mPipe_rData_id <= mBusAxi_aw_s2mPipe_payload_id;
      mBusAxi_aw_s2mPipe_rData_len <= mBusAxi_aw_s2mPipe_payload_len;
      mBusAxi_aw_s2mPipe_rData_size <= mBusAxi_aw_s2mPipe_payload_size;
      mBusAxi_aw_s2mPipe_rData_burst <= mBusAxi_aw_s2mPipe_payload_burst;
      mBusAxi_aw_s2mPipe_rData_allStrb <= mBusAxi_aw_s2mPipe_payload_allStrb;
    end
    if(mBusAxi_w_ready) begin
      mBusAxi_w_rData_data <= mBusAxi_w_payload_data;
      mBusAxi_w_rData_strb <= mBusAxi_w_payload_strb;
      mBusAxi_w_rData_last <= mBusAxi_w_payload_last;
    end
    if(mBusAxi_w_s2mPipe_ready) begin
      mBusAxi_w_s2mPipe_rData_data <= mBusAxi_w_s2mPipe_payload_data;
      mBusAxi_w_s2mPipe_rData_strb <= mBusAxi_w_s2mPipe_payload_strb;
      mBusAxi_w_s2mPipe_rData_last <= mBusAxi_w_s2mPipe_payload_last;
    end
    if(mBus_bready) begin
      mBus_b_rData_id <= mBus_bid;
      mBus_b_rData_resp <= mBus_bresp;
    end
    if(mBus_b_s2mPipe_ready) begin
      mBus_b_s2mPipe_rData_id <= mBus_b_s2mPipe_payload_id;
      mBus_b_s2mPipe_rData_resp <= mBus_b_s2mPipe_payload_resp;
    end
    if(mBusAxi_ar_ready) begin
      mBusAxi_ar_rData_addr <= mBusAxi_ar_payload_addr;
      mBusAxi_ar_rData_id <= mBusAxi_ar_payload_id;
      mBusAxi_ar_rData_len <= mBusAxi_ar_payload_len;
      mBusAxi_ar_rData_size <= mBusAxi_ar_payload_size;
      mBusAxi_ar_rData_burst <= mBusAxi_ar_payload_burst;
    end
    if(mBusAxi_ar_s2mPipe_ready) begin
      mBusAxi_ar_s2mPipe_rData_addr <= mBusAxi_ar_s2mPipe_payload_addr;
      mBusAxi_ar_s2mPipe_rData_id <= mBusAxi_ar_s2mPipe_payload_id;
      mBusAxi_ar_s2mPipe_rData_len <= mBusAxi_ar_s2mPipe_payload_len;
      mBusAxi_ar_s2mPipe_rData_size <= mBusAxi_ar_s2mPipe_payload_size;
      mBusAxi_ar_s2mPipe_rData_burst <= mBusAxi_ar_s2mPipe_payload_burst;
    end
    if(mBus_rready) begin
      mBus_r_rData_data <= mBus_rdata;
      mBus_r_rData_id <= mBus_rid;
      mBus_r_rData_resp <= mBus_rresp;
      mBus_r_rData_last <= mBus_rlast;
    end
    if(mBus_r_s2mPipe_ready) begin
      mBus_r_s2mPipe_rData_data <= mBus_r_s2mPipe_payload_data;
      mBus_r_s2mPipe_rData_id <= mBus_r_s2mPipe_payload_id;
      mBus_r_s2mPipe_rData_resp <= mBus_r_s2mPipe_payload_resp;
      mBus_r_s2mPipe_rData_last <= mBus_r_s2mPipe_payload_last;
    end
    debugIn_delay_1 <= debugIn;
    debug <= debugIn_delay_1;
  end

  always @(posedge litex_clk or posedge cpuResetCtrl_fiber_aggregator_reset) begin
    if(cpuResetCtrl_fiber_aggregator_reset) begin
      cpuResetCtrl_fiber_holder_counter <= 7'h0;
    end else begin
      if(when_CrossClock_l341) begin
        cpuResetCtrl_fiber_holder_counter <= (cpuResetCtrl_fiber_holder_counter + 7'h01);
      end
    end
  end

  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      vexiis_0_dBus_bus_a_rValid <= 1'b0;
      vexiis_0_dBus_noDecoder_toDown_d_rValid <= 1'b0;
      vexiis_0_iBus_bus_a_rValid <= 1'b0;
      vexiis_0_iBus_bus_a_halfPipe_rValid <= 1'b0;
      vexiis_0_iBus_noDecoder_toDown_d_rValid <= 1'b0;
      vexiis_0_lsuL1Bus_bus_a_rValidN <= 1'b1;
      vexiis_0_lsuL1Bus_bus_a_s2mPipe_rValid <= 1'b0;
      vexiis_0_lsuL1Bus_noDecoder_toDown_d_rValid <= 1'b0;
      vexiis_0_dBus_to_ioBus_down_bus_a_rValid <= 1'b0;
      mBusAxi_aw_rValidN <= 1'b1;
      mBusAxi_aw_s2mPipe_rValid <= 1'b0;
      mBusAxi_w_rValidN <= 1'b1;
      mBusAxi_w_s2mPipe_rValid <= 1'b0;
      mBus_b_rValidN <= 1'b1;
      mBus_b_s2mPipe_rValid <= 1'b0;
      mBusAxi_ar_rValidN <= 1'b1;
      mBusAxi_ar_s2mPipe_rValid <= 1'b0;
      mBus_r_rValidN <= 1'b1;
      mBus_r_s2mPipe_rValid <= 1'b0;
    end else begin
      if(vexiis_0_dBus_bus_a_valid) begin
        vexiis_0_dBus_bus_a_rValid <= 1'b1;
      end
      if(vexiis_0_dBus_bus_a_halfPipe_fire) begin
        vexiis_0_dBus_bus_a_rValid <= 1'b0;
      end
      if(vexiis_0_dBus_noDecoder_toDown_d_ready) begin
        vexiis_0_dBus_noDecoder_toDown_d_rValid <= vexiis_0_dBus_noDecoder_toDown_d_valid;
      end
      if(vexiis_0_iBus_bus_a_valid) begin
        vexiis_0_iBus_bus_a_rValid <= 1'b1;
      end
      if(vexiis_0_iBus_bus_a_halfPipe_fire) begin
        vexiis_0_iBus_bus_a_rValid <= 1'b0;
      end
      if(vexiis_0_iBus_bus_a_halfPipe_valid) begin
        vexiis_0_iBus_bus_a_halfPipe_rValid <= 1'b1;
      end
      if(vexiis_0_iBus_bus_a_halfPipe_halfPipe_fire) begin
        vexiis_0_iBus_bus_a_halfPipe_rValid <= 1'b0;
      end
      if(vexiis_0_iBus_noDecoder_toDown_d_ready) begin
        vexiis_0_iBus_noDecoder_toDown_d_rValid <= vexiis_0_iBus_noDecoder_toDown_d_valid;
      end
      if(vexiis_0_lsuL1Bus_bus_a_valid) begin
        vexiis_0_lsuL1Bus_bus_a_rValidN <= 1'b0;
      end
      if(vexiis_0_lsuL1Bus_bus_a_s2mPipe_ready) begin
        vexiis_0_lsuL1Bus_bus_a_rValidN <= 1'b1;
      end
      if(vexiis_0_lsuL1Bus_bus_a_s2mPipe_ready) begin
        vexiis_0_lsuL1Bus_bus_a_s2mPipe_rValid <= vexiis_0_lsuL1Bus_bus_a_s2mPipe_valid;
      end
      if(vexiis_0_lsuL1Bus_noDecoder_toDown_d_ready) begin
        vexiis_0_lsuL1Bus_noDecoder_toDown_d_rValid <= vexiis_0_lsuL1Bus_noDecoder_toDown_d_valid;
      end
      if(vexiis_0_dBus_to_ioBus_down_bus_a_valid) begin
        vexiis_0_dBus_to_ioBus_down_bus_a_rValid <= 1'b1;
      end
      if(vexiis_0_dBus_to_ioBus_down_bus_a_halfPipe_fire) begin
        vexiis_0_dBus_to_ioBus_down_bus_a_rValid <= 1'b0;
      end
      if(mBusAxi_aw_valid) begin
        mBusAxi_aw_rValidN <= 1'b0;
      end
      if(mBusAxi_aw_s2mPipe_ready) begin
        mBusAxi_aw_rValidN <= 1'b1;
      end
      if(mBusAxi_aw_s2mPipe_ready) begin
        mBusAxi_aw_s2mPipe_rValid <= mBusAxi_aw_s2mPipe_valid;
      end
      if(mBusAxi_w_valid) begin
        mBusAxi_w_rValidN <= 1'b0;
      end
      if(mBusAxi_w_s2mPipe_ready) begin
        mBusAxi_w_rValidN <= 1'b1;
      end
      if(mBusAxi_w_s2mPipe_ready) begin
        mBusAxi_w_s2mPipe_rValid <= mBusAxi_w_s2mPipe_valid;
      end
      if(mBus_bvalid) begin
        mBus_b_rValidN <= 1'b0;
      end
      if(mBus_b_s2mPipe_ready) begin
        mBus_b_rValidN <= 1'b1;
      end
      if(mBus_b_s2mPipe_ready) begin
        mBus_b_s2mPipe_rValid <= mBus_b_s2mPipe_valid;
      end
      if(mBusAxi_ar_valid) begin
        mBusAxi_ar_rValidN <= 1'b0;
      end
      if(mBusAxi_ar_s2mPipe_ready) begin
        mBusAxi_ar_rValidN <= 1'b1;
      end
      if(mBusAxi_ar_s2mPipe_ready) begin
        mBusAxi_ar_s2mPipe_rValid <= mBusAxi_ar_s2mPipe_valid;
      end
      if(mBus_rvalid) begin
        mBus_r_rValidN <= 1'b0;
      end
      if(mBus_r_s2mPipe_ready) begin
        mBus_r_rValidN <= 1'b1;
      end
      if(mBus_r_s2mPipe_ready) begin
        mBus_r_s2mPipe_rValid <= mBus_r_s2mPipe_valid;
      end
    end
  end

  always @(posedge litex_clk or posedge litex_reset) begin
    if(litex_reset) begin
      peripheral_bus_bus_a_rValid <= 1'b0;
      io_up_d_rValid <= 1'b0;
      peripheral_toAxiLite4_down_aw_rValid <= 1'b0;
      peripheral_toAxiLite4_down_w_rValid <= 1'b0;
      pBus_b_rValid <= 1'b0;
      peripheral_toAxiLite4_down_ar_rValid <= 1'b0;
      pBus_r_rValid <= 1'b0;
    end else begin
      if(peripheral_bus_bus_a_valid) begin
        peripheral_bus_bus_a_rValid <= 1'b1;
      end
      if(peripheral_bus_bus_a_halfPipe_fire) begin
        peripheral_bus_bus_a_rValid <= 1'b0;
      end
      if(peripheral_bus_decoder_core_io_up_d_valid) begin
        io_up_d_rValid <= 1'b1;
      end
      if(io_up_d_halfPipe_fire) begin
        io_up_d_rValid <= 1'b0;
      end
      if(peripheral_toAxiLite4_down_aw_valid) begin
        peripheral_toAxiLite4_down_aw_rValid <= 1'b1;
      end
      if(peripheral_toAxiLite4_down_aw_halfPipe_fire) begin
        peripheral_toAxiLite4_down_aw_rValid <= 1'b0;
      end
      if(peripheral_toAxiLite4_down_w_valid) begin
        peripheral_toAxiLite4_down_w_rValid <= 1'b1;
      end
      if(peripheral_toAxiLite4_down_w_halfPipe_fire) begin
        peripheral_toAxiLite4_down_w_rValid <= 1'b0;
      end
      if(pBus_bvalid) begin
        pBus_b_rValid <= 1'b1;
      end
      if(pBus_b_halfPipe_fire) begin
        pBus_b_rValid <= 1'b0;
      end
      if(peripheral_toAxiLite4_down_ar_valid) begin
        peripheral_toAxiLite4_down_ar_rValid <= 1'b1;
      end
      if(peripheral_toAxiLite4_down_ar_halfPipe_fire) begin
        peripheral_toAxiLite4_down_ar_rValid <= 1'b0;
      end
      if(pBus_rvalid) begin
        pBus_r_rValid <= 1'b1;
      end
      if(pBus_r_halfPipe_fire) begin
        pBus_r_rValid <= 1'b0;
      end
    end
  end

  always @(posedge litex_clk) begin
    if(peripheral_bus_bus_a_ready) begin
      peripheral_bus_bus_a_rData_opcode <= peripheral_bus_bus_a_payload_opcode;
      peripheral_bus_bus_a_rData_param <= peripheral_bus_bus_a_payload_param;
      peripheral_bus_bus_a_rData_source <= peripheral_bus_bus_a_payload_source;
      peripheral_bus_bus_a_rData_address <= peripheral_bus_bus_a_payload_address;
      peripheral_bus_bus_a_rData_size <= peripheral_bus_bus_a_payload_size;
      peripheral_bus_bus_a_rData_mask <= peripheral_bus_bus_a_payload_mask;
      peripheral_bus_bus_a_rData_data <= peripheral_bus_bus_a_payload_data;
      peripheral_bus_bus_a_rData_corrupt <= peripheral_bus_bus_a_payload_corrupt;
    end
    if(peripheral_bus_decoder_core_io_up_d_ready) begin
      io_up_d_rData_opcode <= peripheral_bus_decoder_core_io_up_d_payload_opcode;
      io_up_d_rData_param <= peripheral_bus_decoder_core_io_up_d_payload_param;
      io_up_d_rData_source <= peripheral_bus_decoder_core_io_up_d_payload_source;
      io_up_d_rData_size <= peripheral_bus_decoder_core_io_up_d_payload_size;
      io_up_d_rData_denied <= peripheral_bus_decoder_core_io_up_d_payload_denied;
      io_up_d_rData_data <= peripheral_bus_decoder_core_io_up_d_payload_data;
      io_up_d_rData_corrupt <= peripheral_bus_decoder_core_io_up_d_payload_corrupt;
    end
    if(peripheral_toAxiLite4_down_aw_ready) begin
      peripheral_toAxiLite4_down_aw_rData_addr <= peripheral_toAxiLite4_down_aw_payload_addr;
      peripheral_toAxiLite4_down_aw_rData_prot <= peripheral_toAxiLite4_down_aw_payload_prot;
    end
    if(peripheral_toAxiLite4_down_w_ready) begin
      peripheral_toAxiLite4_down_w_rData_data <= peripheral_toAxiLite4_down_w_payload_data;
      peripheral_toAxiLite4_down_w_rData_strb <= peripheral_toAxiLite4_down_w_payload_strb;
    end
    if(pBus_bready) begin
      pBus_b_rData_resp <= pBus_bresp;
    end
    if(peripheral_toAxiLite4_down_ar_ready) begin
      peripheral_toAxiLite4_down_ar_rData_addr <= peripheral_toAxiLite4_down_ar_payload_addr;
      peripheral_toAxiLite4_down_ar_rData_prot <= peripheral_toAxiLite4_down_ar_payload_prot;
    end
    if(pBus_rready) begin
      pBus_r_rData_data <= pBus_rdata;
      pBus_r_rData_resp <= pBus_rresp;
    end
  end


endmodule

module Decoder_1 (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [2:0]    io_up_a_payload_source,
  input  wire [31:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [3:0]    io_up_a_payload_mask,
  input  wire [31:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [2:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [31:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_downs_0_a_valid,
  input  wire          io_downs_0_a_ready,
  output wire [2:0]    io_downs_0_a_payload_opcode,
  output wire [2:0]    io_downs_0_a_payload_param,
  output wire [2:0]    io_downs_0_a_payload_source,
  output wire [15:0]   io_downs_0_a_payload_address,
  output wire [2:0]    io_downs_0_a_payload_size,
  output wire [3:0]    io_downs_0_a_payload_mask,
  output wire [31:0]   io_downs_0_a_payload_data,
  output wire          io_downs_0_a_payload_corrupt,
  input  wire          io_downs_0_d_valid,
  output wire          io_downs_0_d_ready,
  input  wire [2:0]    io_downs_0_d_payload_opcode,
  input  wire [2:0]    io_downs_0_d_payload_param,
  input  wire [2:0]    io_downs_0_d_payload_source,
  input  wire [2:0]    io_downs_0_d_payload_size,
  input  wire          io_downs_0_d_payload_denied,
  input  wire [31:0]   io_downs_0_d_payload_data,
  input  wire          io_downs_0_d_payload_corrupt,
  output wire          io_downs_1_a_valid,
  input  wire          io_downs_1_a_ready,
  output wire [2:0]    io_downs_1_a_payload_opcode,
  output wire [2:0]    io_downs_1_a_payload_param,
  output wire [2:0]    io_downs_1_a_payload_source,
  output wire [21:0]   io_downs_1_a_payload_address,
  output wire [1:0]    io_downs_1_a_payload_size,
  output wire [3:0]    io_downs_1_a_payload_mask,
  output wire [31:0]   io_downs_1_a_payload_data,
  output wire          io_downs_1_a_payload_corrupt,
  input  wire          io_downs_1_d_valid,
  output wire          io_downs_1_d_ready,
  input  wire [2:0]    io_downs_1_d_payload_opcode,
  input  wire [2:0]    io_downs_1_d_payload_param,
  input  wire [2:0]    io_downs_1_d_payload_source,
  input  wire [1:0]    io_downs_1_d_payload_size,
  input  wire          io_downs_1_d_payload_denied,
  input  wire [31:0]   io_downs_1_d_payload_data,
  input  wire          io_downs_1_d_payload_corrupt,
  output wire          io_downs_2_a_valid,
  input  wire          io_downs_2_a_ready,
  output wire [2:0]    io_downs_2_a_payload_opcode,
  output wire [2:0]    io_downs_2_a_payload_param,
  output wire [2:0]    io_downs_2_a_payload_source,
  output wire [31:0]   io_downs_2_a_payload_address,
  output wire [2:0]    io_downs_2_a_payload_size,
  output wire [3:0]    io_downs_2_a_payload_mask,
  output wire [31:0]   io_downs_2_a_payload_data,
  output wire          io_downs_2_a_payload_corrupt,
  input  wire          io_downs_2_d_valid,
  output wire          io_downs_2_d_ready,
  input  wire [2:0]    io_downs_2_d_payload_opcode,
  input  wire [2:0]    io_downs_2_d_payload_param,
  input  wire [2:0]    io_downs_2_d_payload_source,
  input  wire [2:0]    io_downs_2_d_payload_size,
  input  wire          io_downs_2_d_payload_denied,
  input  wire [31:0]   io_downs_2_d_payload_data,
  input  wire          io_downs_2_d_payload_corrupt,
  input  wire          litex_clk,
  input  wire          litex_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire       [2:0]    d_arbiter_io_inputs_1_payload_size;
  wire                d_arbiter_io_inputs_0_ready;
  wire                d_arbiter_io_inputs_1_ready;
  wire                d_arbiter_io_inputs_2_ready;
  wire                d_arbiter_io_output_valid;
  wire       [2:0]    d_arbiter_io_output_payload_opcode;
  wire       [2:0]    d_arbiter_io_output_payload_param;
  wire       [2:0]    d_arbiter_io_output_payload_source;
  wire       [2:0]    d_arbiter_io_output_payload_size;
  wire                d_arbiter_io_output_payload_denied;
  wire       [31:0]   d_arbiter_io_output_payload_data;
  wire                d_arbiter_io_output_payload_corrupt;
  wire       [1:0]    d_arbiter_io_chosen;
  wire       [2:0]    d_arbiter_io_chosenOH;
  wire       [0:0]    _zz_a_logic_0_hit;
  wire       [31:0]   _zz_downs_0_a_payload_address;
  wire       [0:0]    _zz_a_logic_1_hit;
  wire       [31:0]   _zz_downs_1_a_payload_address;
  wire       [0:0]    _zz_a_logic_2_hit;
  reg        [1:0]    _zz_1;
  wire       [2:0]    _zz_2;
  wire                downs_0_a_valid;
  wire                downs_0_a_ready;
  wire       [2:0]    downs_0_a_payload_opcode;
  wire       [2:0]    downs_0_a_payload_param;
  wire       [2:0]    downs_0_a_payload_source;
  wire       [15:0]   downs_0_a_payload_address;
  wire       [2:0]    downs_0_a_payload_size;
  wire       [3:0]    downs_0_a_payload_mask;
  wire       [31:0]   downs_0_a_payload_data;
  wire                downs_0_a_payload_corrupt;
  wire                downs_0_d_valid;
  wire                downs_0_d_ready;
  wire       [2:0]    downs_0_d_payload_opcode;
  wire       [2:0]    downs_0_d_payload_param;
  wire       [2:0]    downs_0_d_payload_source;
  wire       [2:0]    downs_0_d_payload_size;
  wire                downs_0_d_payload_denied;
  wire       [31:0]   downs_0_d_payload_data;
  wire                downs_0_d_payload_corrupt;
  wire                downs_1_a_valid;
  wire                downs_1_a_ready;
  wire       [2:0]    downs_1_a_payload_opcode;
  wire       [2:0]    downs_1_a_payload_param;
  wire       [2:0]    downs_1_a_payload_source;
  wire       [21:0]   downs_1_a_payload_address;
  wire       [1:0]    downs_1_a_payload_size;
  wire       [3:0]    downs_1_a_payload_mask;
  wire       [31:0]   downs_1_a_payload_data;
  wire                downs_1_a_payload_corrupt;
  wire                downs_1_d_valid;
  wire                downs_1_d_ready;
  wire       [2:0]    downs_1_d_payload_opcode;
  wire       [2:0]    downs_1_d_payload_param;
  wire       [2:0]    downs_1_d_payload_source;
  wire       [1:0]    downs_1_d_payload_size;
  wire                downs_1_d_payload_denied;
  wire       [31:0]   downs_1_d_payload_data;
  wire                downs_1_d_payload_corrupt;
  wire                downs_2_a_valid;
  wire                downs_2_a_ready;
  wire       [2:0]    downs_2_a_payload_opcode;
  wire       [2:0]    downs_2_a_payload_param;
  wire       [2:0]    downs_2_a_payload_source;
  wire       [31:0]   downs_2_a_payload_address;
  wire       [2:0]    downs_2_a_payload_size;
  wire       [3:0]    downs_2_a_payload_mask;
  wire       [31:0]   downs_2_a_payload_data;
  wire                downs_2_a_payload_corrupt;
  wire                downs_2_d_valid;
  wire                downs_2_d_ready;
  wire       [2:0]    downs_2_d_payload_opcode;
  wire       [2:0]    downs_2_d_payload_param;
  wire       [2:0]    downs_2_d_payload_source;
  wire       [2:0]    downs_2_d_payload_size;
  wire                downs_2_d_payload_denied;
  wire       [31:0]   downs_2_d_payload_data;
  wire                downs_2_d_payload_corrupt;
  wire       [34:0]   a_key;
  wire                a_logic_0_hit;
  wire                a_logic_1_hit;
  wire                a_logic_2_hit;
  wire                a_miss;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] io_downs_0_a_payload_opcode_string;
  reg [119:0] io_downs_0_d_payload_opcode_string;
  reg [127:0] io_downs_1_a_payload_opcode_string;
  reg [119:0] io_downs_1_d_payload_opcode_string;
  reg [127:0] io_downs_2_a_payload_opcode_string;
  reg [119:0] io_downs_2_d_payload_opcode_string;
  reg [127:0] downs_0_a_payload_opcode_string;
  reg [119:0] downs_0_d_payload_opcode_string;
  reg [127:0] downs_1_a_payload_opcode_string;
  reg [119:0] downs_1_d_payload_opcode_string;
  reg [127:0] downs_2_a_payload_opcode_string;
  reg [119:0] downs_2_d_payload_opcode_string;
  `endif


  assign _zz_a_logic_0_hit = (|((a_key & 35'h001810000) == 35'h000010000));
  assign _zz_downs_0_a_payload_address = (io_up_a_payload_address - 32'hf0010000);
  assign _zz_a_logic_1_hit = (|((a_key & 35'h001800000) == 35'h000800000));
  assign _zz_downs_1_a_payload_address = (io_up_a_payload_address - 32'hf0c00000);
  assign _zz_a_logic_2_hit = (|{((a_key & 35'h080000000) == 35'h0),((a_key & 35'h000810000) == 35'h0)});
  assign _zz_2 = {io_downs_2_a_valid,{io_downs_1_a_valid,io_downs_0_a_valid}};
  StreamArbiter_9 d_arbiter (
    .io_inputs_0_valid           (downs_0_d_valid                        ), //i
    .io_inputs_0_ready           (d_arbiter_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_opcode  (downs_0_d_payload_opcode[2:0]          ), //i
    .io_inputs_0_payload_param   (downs_0_d_payload_param[2:0]           ), //i
    .io_inputs_0_payload_source  (downs_0_d_payload_source[2:0]          ), //i
    .io_inputs_0_payload_size    (downs_0_d_payload_size[2:0]            ), //i
    .io_inputs_0_payload_denied  (downs_0_d_payload_denied               ), //i
    .io_inputs_0_payload_data    (downs_0_d_payload_data[31:0]           ), //i
    .io_inputs_0_payload_corrupt (downs_0_d_payload_corrupt              ), //i
    .io_inputs_1_valid           (downs_1_d_valid                        ), //i
    .io_inputs_1_ready           (d_arbiter_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_opcode  (downs_1_d_payload_opcode[2:0]          ), //i
    .io_inputs_1_payload_param   (downs_1_d_payload_param[2:0]           ), //i
    .io_inputs_1_payload_source  (downs_1_d_payload_source[2:0]          ), //i
    .io_inputs_1_payload_size    (d_arbiter_io_inputs_1_payload_size[2:0]), //i
    .io_inputs_1_payload_denied  (downs_1_d_payload_denied               ), //i
    .io_inputs_1_payload_data    (downs_1_d_payload_data[31:0]           ), //i
    .io_inputs_1_payload_corrupt (downs_1_d_payload_corrupt              ), //i
    .io_inputs_2_valid           (downs_2_d_valid                        ), //i
    .io_inputs_2_ready           (d_arbiter_io_inputs_2_ready            ), //o
    .io_inputs_2_payload_opcode  (downs_2_d_payload_opcode[2:0]          ), //i
    .io_inputs_2_payload_param   (downs_2_d_payload_param[2:0]           ), //i
    .io_inputs_2_payload_source  (downs_2_d_payload_source[2:0]          ), //i
    .io_inputs_2_payload_size    (downs_2_d_payload_size[2:0]            ), //i
    .io_inputs_2_payload_denied  (downs_2_d_payload_denied               ), //i
    .io_inputs_2_payload_data    (downs_2_d_payload_data[31:0]           ), //i
    .io_inputs_2_payload_corrupt (downs_2_d_payload_corrupt              ), //i
    .io_output_valid             (d_arbiter_io_output_valid              ), //o
    .io_output_ready             (io_up_d_ready                          ), //i
    .io_output_payload_opcode    (d_arbiter_io_output_payload_opcode[2:0]), //o
    .io_output_payload_param     (d_arbiter_io_output_payload_param[2:0] ), //o
    .io_output_payload_source    (d_arbiter_io_output_payload_source[2:0]), //o
    .io_output_payload_size      (d_arbiter_io_output_payload_size[2:0]  ), //o
    .io_output_payload_denied    (d_arbiter_io_output_payload_denied     ), //o
    .io_output_payload_data      (d_arbiter_io_output_payload_data[31:0] ), //o
    .io_output_payload_corrupt   (d_arbiter_io_output_payload_corrupt    ), //o
    .io_chosen                   (d_arbiter_io_chosen[1:0]               ), //o
    .io_chosenOH                 (d_arbiter_io_chosenOH[2:0]             ), //o
    .litex_clk                   (litex_clk                              ), //i
    .litex_reset                 (litex_reset                            )  //i
  );
  always @(*) begin
    case(_zz_2)
      3'b000 : _zz_1 = 2'b00;
      3'b001 : _zz_1 = 2'b01;
      3'b010 : _zz_1 = 2'b01;
      3'b011 : _zz_1 = 2'b10;
      3'b100 : _zz_1 = 2'b01;
      3'b101 : _zz_1 = 2'b10;
      3'b110 : _zz_1 = 2'b10;
      default : _zz_1 = 2'b11;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_0_a_payload_opcode)
      A_PUT_FULL_DATA : io_downs_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_downs_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_downs_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_downs_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_downs_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_downs_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_0_d_payload_opcode)
      D_ACCESS_ACK : io_downs_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_downs_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_downs_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_downs_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_downs_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_downs_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_1_a_payload_opcode)
      A_PUT_FULL_DATA : io_downs_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_downs_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_downs_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_downs_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_downs_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_downs_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_1_d_payload_opcode)
      D_ACCESS_ACK : io_downs_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_downs_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_downs_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_downs_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_downs_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_downs_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_2_a_payload_opcode)
      A_PUT_FULL_DATA : io_downs_2_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_downs_2_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_downs_2_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_downs_2_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_downs_2_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_downs_2_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_2_d_payload_opcode)
      D_ACCESS_ACK : io_downs_2_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_downs_2_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_downs_2_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_downs_2_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_downs_2_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_downs_2_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downs_0_a_payload_opcode)
      A_PUT_FULL_DATA : downs_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downs_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downs_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downs_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downs_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : downs_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(downs_0_d_payload_opcode)
      D_ACCESS_ACK : downs_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : downs_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : downs_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : downs_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : downs_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : downs_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downs_1_a_payload_opcode)
      A_PUT_FULL_DATA : downs_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downs_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downs_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downs_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downs_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : downs_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(downs_1_d_payload_opcode)
      D_ACCESS_ACK : downs_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : downs_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : downs_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : downs_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : downs_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : downs_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downs_2_a_payload_opcode)
      A_PUT_FULL_DATA : downs_2_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downs_2_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downs_2_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downs_2_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downs_2_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : downs_2_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(downs_2_d_payload_opcode)
      D_ACCESS_ACK : downs_2_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : downs_2_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : downs_2_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : downs_2_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : downs_2_d_payload_opcode_string = "RELEASE_ACK    ";
      default : downs_2_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign io_downs_0_a_valid = downs_0_a_valid;
  assign downs_0_a_ready = io_downs_0_a_ready;
  assign io_downs_0_a_payload_opcode = downs_0_a_payload_opcode;
  assign io_downs_0_a_payload_param = downs_0_a_payload_param;
  assign io_downs_0_a_payload_source = downs_0_a_payload_source;
  assign io_downs_0_a_payload_address = downs_0_a_payload_address;
  assign io_downs_0_a_payload_size = downs_0_a_payload_size;
  assign io_downs_0_a_payload_mask = downs_0_a_payload_mask;
  assign io_downs_0_a_payload_data = downs_0_a_payload_data;
  assign io_downs_0_a_payload_corrupt = downs_0_a_payload_corrupt;
  assign downs_0_d_valid = io_downs_0_d_valid;
  assign io_downs_0_d_ready = downs_0_d_ready;
  assign downs_0_d_payload_opcode = io_downs_0_d_payload_opcode;
  assign downs_0_d_payload_param = io_downs_0_d_payload_param;
  assign downs_0_d_payload_source = io_downs_0_d_payload_source;
  assign downs_0_d_payload_size = io_downs_0_d_payload_size;
  assign downs_0_d_payload_denied = io_downs_0_d_payload_denied;
  assign downs_0_d_payload_data = io_downs_0_d_payload_data;
  assign downs_0_d_payload_corrupt = io_downs_0_d_payload_corrupt;
  assign io_downs_1_a_valid = downs_1_a_valid;
  assign downs_1_a_ready = io_downs_1_a_ready;
  assign io_downs_1_a_payload_opcode = downs_1_a_payload_opcode;
  assign io_downs_1_a_payload_param = downs_1_a_payload_param;
  assign io_downs_1_a_payload_source = downs_1_a_payload_source;
  assign io_downs_1_a_payload_address = downs_1_a_payload_address;
  assign io_downs_1_a_payload_size = downs_1_a_payload_size;
  assign io_downs_1_a_payload_mask = downs_1_a_payload_mask;
  assign io_downs_1_a_payload_data = downs_1_a_payload_data;
  assign io_downs_1_a_payload_corrupt = downs_1_a_payload_corrupt;
  assign downs_1_d_valid = io_downs_1_d_valid;
  assign io_downs_1_d_ready = downs_1_d_ready;
  assign downs_1_d_payload_opcode = io_downs_1_d_payload_opcode;
  assign downs_1_d_payload_param = io_downs_1_d_payload_param;
  assign downs_1_d_payload_source = io_downs_1_d_payload_source;
  assign downs_1_d_payload_size = io_downs_1_d_payload_size;
  assign downs_1_d_payload_denied = io_downs_1_d_payload_denied;
  assign downs_1_d_payload_data = io_downs_1_d_payload_data;
  assign downs_1_d_payload_corrupt = io_downs_1_d_payload_corrupt;
  assign io_downs_2_a_valid = downs_2_a_valid;
  assign downs_2_a_ready = io_downs_2_a_ready;
  assign io_downs_2_a_payload_opcode = downs_2_a_payload_opcode;
  assign io_downs_2_a_payload_param = downs_2_a_payload_param;
  assign io_downs_2_a_payload_source = downs_2_a_payload_source;
  assign io_downs_2_a_payload_address = downs_2_a_payload_address;
  assign io_downs_2_a_payload_size = downs_2_a_payload_size;
  assign io_downs_2_a_payload_mask = downs_2_a_payload_mask;
  assign io_downs_2_a_payload_data = downs_2_a_payload_data;
  assign io_downs_2_a_payload_corrupt = downs_2_a_payload_corrupt;
  assign downs_2_d_valid = io_downs_2_d_valid;
  assign io_downs_2_d_ready = downs_2_d_ready;
  assign downs_2_d_payload_opcode = io_downs_2_d_payload_opcode;
  assign downs_2_d_payload_param = io_downs_2_d_payload_param;
  assign downs_2_d_payload_source = io_downs_2_d_payload_source;
  assign downs_2_d_payload_size = io_downs_2_d_payload_size;
  assign downs_2_d_payload_denied = io_downs_2_d_payload_denied;
  assign downs_2_d_payload_data = io_downs_2_d_payload_data;
  assign downs_2_d_payload_corrupt = io_downs_2_d_payload_corrupt;
  assign a_key = {io_up_a_payload_opcode,io_up_a_payload_address};
  assign a_logic_0_hit = _zz_a_logic_0_hit[0];
  assign downs_0_a_valid = (io_up_a_valid && a_logic_0_hit);
  assign downs_0_a_payload_opcode = io_up_a_payload_opcode;
  assign downs_0_a_payload_param = io_up_a_payload_param;
  assign downs_0_a_payload_source = io_up_a_payload_source;
  assign downs_0_a_payload_mask = io_up_a_payload_mask;
  assign downs_0_a_payload_data = io_up_a_payload_data;
  assign downs_0_a_payload_corrupt = io_up_a_payload_corrupt;
  assign downs_0_a_payload_address = _zz_downs_0_a_payload_address[15:0];
  assign downs_0_a_payload_size = io_up_a_payload_size;
  assign a_logic_1_hit = _zz_a_logic_1_hit[0];
  assign downs_1_a_valid = (io_up_a_valid && a_logic_1_hit);
  assign downs_1_a_payload_opcode = io_up_a_payload_opcode;
  assign downs_1_a_payload_param = io_up_a_payload_param;
  assign downs_1_a_payload_source = io_up_a_payload_source;
  assign downs_1_a_payload_mask = io_up_a_payload_mask;
  assign downs_1_a_payload_data = io_up_a_payload_data;
  assign downs_1_a_payload_corrupt = io_up_a_payload_corrupt;
  assign downs_1_a_payload_address = _zz_downs_1_a_payload_address[21:0];
  assign downs_1_a_payload_size = io_up_a_payload_size[1:0];
  assign a_logic_2_hit = _zz_a_logic_2_hit[0];
  assign downs_2_a_valid = (io_up_a_valid && a_logic_2_hit);
  assign downs_2_a_payload_opcode = io_up_a_payload_opcode;
  assign downs_2_a_payload_param = io_up_a_payload_param;
  assign downs_2_a_payload_source = io_up_a_payload_source;
  assign downs_2_a_payload_mask = io_up_a_payload_mask;
  assign downs_2_a_payload_data = io_up_a_payload_data;
  assign downs_2_a_payload_corrupt = io_up_a_payload_corrupt;
  assign downs_2_a_payload_address = io_up_a_payload_address;
  assign downs_2_a_payload_size = io_up_a_payload_size;
  assign io_up_a_ready = (|{(downs_2_a_ready && a_logic_2_hit),{(downs_1_a_ready && a_logic_1_hit),(downs_0_a_ready && a_logic_0_hit)}});
  assign a_miss = (! (|{a_logic_2_hit,{a_logic_1_hit,a_logic_0_hit}}));
  assign downs_0_d_ready = d_arbiter_io_inputs_0_ready;
  assign downs_1_d_ready = d_arbiter_io_inputs_1_ready;
  assign d_arbiter_io_inputs_1_payload_size = {1'd0, downs_1_d_payload_size};
  assign downs_2_d_ready = d_arbiter_io_inputs_2_ready;
  assign io_up_d_valid = d_arbiter_io_output_valid;
  assign io_up_d_payload_opcode = d_arbiter_io_output_payload_opcode;
  assign io_up_d_payload_param = d_arbiter_io_output_payload_param;
  assign io_up_d_payload_source = d_arbiter_io_output_payload_source;
  assign io_up_d_payload_size = d_arbiter_io_output_payload_size;
  assign io_up_d_payload_denied = d_arbiter_io_output_payload_denied;
  assign io_up_d_payload_data = d_arbiter_io_output_payload_data;
  assign io_up_d_payload_corrupt = d_arbiter_io_output_payload_corrupt;
  always @(posedge litex_clk or posedge litex_reset) begin
    if(litex_reset) begin
    end else begin
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (io_up_a_valid && a_miss))); // Decoder.scala:L106
        `else
          if(!(! (io_up_a_valid && a_miss))) begin
            $display("FAILURE Tilelink decoder miss ???"); // Decoder.scala:L106
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (io_up_a_valid && (_zz_1 != 2'b01)))); // Decoder.scala:L107
        `else
          if(!(! (io_up_a_valid && (_zz_1 != 2'b01)))) begin
            $display("FAILURE Tilelink decoder miss ???"); // Decoder.scala:L107
            $finish;
          end
        `endif
      `endif
    end
  end


endmodule

module WidthAdapter_1 (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [1:0]    io_up_a_payload_source,
  input  wire [31:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [7:0]    io_up_a_payload_mask,
  input  wire [63:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [1:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [63:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_down_a_valid,
  input  wire          io_down_a_ready,
  output wire [2:0]    io_down_a_payload_opcode,
  output wire [2:0]    io_down_a_payload_param,
  output wire [1:0]    io_down_a_payload_source,
  output reg  [31:0]   io_down_a_payload_address,
  output wire [2:0]    io_down_a_payload_size,
  output wire [3:0]    io_down_a_payload_mask,
  output wire [31:0]   io_down_a_payload_data,
  output wire          io_down_a_payload_corrupt,
  input  wire          io_down_d_valid,
  output wire          io_down_d_ready,
  input  wire [2:0]    io_down_d_payload_opcode,
  input  wire [2:0]    io_down_d_payload_param,
  input  wire [1:0]    io_down_d_payload_source,
  input  wire [2:0]    io_down_d_payload_size,
  input  wire          io_down_d_payload_denied,
  input  wire [31:0]   io_down_d_payload_data,
  input  wire          io_down_d_payload_corrupt,
  input  wire          litex_clk,
  input  wire          litex_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  reg        [3:0]    _zz_downsize_a_ctrl_burstLast;
  reg        [31:0]   _zz_io_down_a_payload_data;
  reg        [3:0]    _zz_io_down_a_payload_mask;
  reg        [3:0]    _zz_downsize_d_ctrl_burstLast;
  reg        [0:0]    downsize_a_ctrl_counter;
  wire       [0:0]    downsize_a_ctrl_sel;
  reg        [3:0]    io_down_a_tracker_beat;
  wire                downsize_a_ctrl_burstLast;
  wire                io_down_a_fire;
  reg        [3:0]    io_down_d_tracker_beat;
  wire                downsize_d_ctrl_burstLast;
  wire                io_down_d_fire;
  wire       [0:0]    downsize_d_sel;
  wire                downsize_d_ctrl_wordLast;
  reg                 downsize_d_ctrl_buffer_valid;
  reg                 downsize_d_ctrl_buffer_first;
  reg        [2:0]    downsize_d_ctrl_buffer_args_opcode;
  reg        [2:0]    downsize_d_ctrl_buffer_args_param;
  reg        [1:0]    downsize_d_ctrl_buffer_args_source;
  reg        [31:0]   downsize_d_ctrl_buffer_args_address;
  reg        [2:0]    downsize_d_ctrl_buffer_args_size;
  reg        [31:0]   downsize_d_ctrl_buffer_data_0;
  reg        [31:0]   downsize_d_ctrl_buffer_data_1;
  reg                 downsize_d_ctrl_buffer_corrupt;
  reg                 downsize_d_ctrl_buffer_denied;
  wire       [0:0]    _zz_when_WidthAdapter_l84;
  wire                when_WidthAdapter_l84;
  wire                when_WidthAdapter_l84_1;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] io_down_a_payload_opcode_string;
  reg [119:0] io_down_d_payload_opcode_string;
  reg [127:0] downsize_d_ctrl_buffer_args_opcode_string;
  `endif


  always @(*) begin
    case(io_down_a_payload_size)
      3'b000 : _zz_downsize_a_ctrl_burstLast = 4'b0000;
      3'b001 : _zz_downsize_a_ctrl_burstLast = 4'b0000;
      3'b010 : _zz_downsize_a_ctrl_burstLast = 4'b0000;
      3'b011 : _zz_downsize_a_ctrl_burstLast = 4'b0001;
      3'b100 : _zz_downsize_a_ctrl_burstLast = 4'b0011;
      3'b101 : _zz_downsize_a_ctrl_burstLast = 4'b0111;
      default : _zz_downsize_a_ctrl_burstLast = 4'b1111;
    endcase
  end

  always @(*) begin
    case(downsize_a_ctrl_sel)
      1'b0 : begin
        _zz_io_down_a_payload_data = io_up_a_payload_data[31 : 0];
        _zz_io_down_a_payload_mask = io_up_a_payload_mask[3 : 0];
      end
      default : begin
        _zz_io_down_a_payload_data = io_up_a_payload_data[63 : 32];
        _zz_io_down_a_payload_mask = io_up_a_payload_mask[7 : 4];
      end
    endcase
  end

  always @(*) begin
    case(io_down_d_payload_size)
      3'b000 : _zz_downsize_d_ctrl_burstLast = 4'b0000;
      3'b001 : _zz_downsize_d_ctrl_burstLast = 4'b0000;
      3'b010 : _zz_downsize_d_ctrl_burstLast = 4'b0000;
      3'b011 : _zz_downsize_d_ctrl_burstLast = 4'b0001;
      3'b100 : _zz_downsize_d_ctrl_burstLast = 4'b0011;
      3'b101 : _zz_downsize_d_ctrl_burstLast = 4'b0111;
      default : _zz_downsize_d_ctrl_burstLast = 4'b1111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_down_a_payload_opcode)
      A_PUT_FULL_DATA : io_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_down_d_payload_opcode)
      D_ACCESS_ACK : io_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downsize_d_ctrl_buffer_args_opcode)
      A_PUT_FULL_DATA : downsize_d_ctrl_buffer_args_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downsize_d_ctrl_buffer_args_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downsize_d_ctrl_buffer_args_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downsize_d_ctrl_buffer_args_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downsize_d_ctrl_buffer_args_opcode_string = "ACQUIRE_PERM    ";
      default : downsize_d_ctrl_buffer_args_opcode_string = "????????????????";
    endcase
  end
  `endif

  assign downsize_a_ctrl_sel = (downsize_a_ctrl_counter + io_up_a_payload_address[2 : 2]);
  assign downsize_a_ctrl_burstLast = ((! ((1'b0 || (A_PUT_FULL_DATA == io_down_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_down_a_payload_opcode))) || (io_down_a_tracker_beat == _zz_downsize_a_ctrl_burstLast));
  assign io_down_a_fire = (io_down_a_valid && io_down_a_ready);
  assign io_down_a_valid = io_up_a_valid;
  assign io_down_a_payload_opcode = io_up_a_payload_opcode;
  assign io_down_a_payload_param = io_up_a_payload_param;
  assign io_down_a_payload_source = io_up_a_payload_source;
  always @(*) begin
    io_down_a_payload_address = io_up_a_payload_address;
    io_down_a_payload_address[2 : 2] = downsize_a_ctrl_sel;
  end

  assign io_down_a_payload_size = io_up_a_payload_size;
  assign io_down_a_payload_corrupt = io_up_a_payload_corrupt;
  assign io_up_a_ready = (io_down_a_ready && ((&downsize_a_ctrl_counter) || downsize_a_ctrl_burstLast));
  assign io_down_a_payload_data = _zz_io_down_a_payload_data;
  assign io_down_a_payload_mask = _zz_io_down_a_payload_mask;
  assign downsize_d_ctrl_burstLast = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_down_d_payload_opcode)) || (D_GRANT_DATA == io_down_d_payload_opcode))) || (io_down_d_tracker_beat == _zz_downsize_d_ctrl_burstLast));
  assign io_down_d_fire = (io_down_d_valid && io_down_d_ready);
  assign downsize_d_sel = io_down_d_tracker_beat[0:0];
  assign downsize_d_ctrl_wordLast = ((&downsize_d_sel) || downsize_d_ctrl_burstLast);
  assign io_up_d_valid = downsize_d_ctrl_buffer_valid;
  assign io_up_d_payload_opcode = downsize_d_ctrl_buffer_args_opcode;
  assign io_up_d_payload_param = downsize_d_ctrl_buffer_args_param;
  assign io_up_d_payload_source = downsize_d_ctrl_buffer_args_source;
  assign io_up_d_payload_size = downsize_d_ctrl_buffer_args_size;
  assign io_up_d_payload_data = {downsize_d_ctrl_buffer_data_1,downsize_d_ctrl_buffer_data_0};
  assign io_up_d_payload_corrupt = downsize_d_ctrl_buffer_corrupt;
  assign io_up_d_payload_denied = downsize_d_ctrl_buffer_denied;
  assign io_down_d_ready = ((! downsize_d_ctrl_buffer_valid) || io_up_d_ready);
  assign _zz_when_WidthAdapter_l84 = (3'b011 <= io_down_d_payload_size);
  assign when_WidthAdapter_l84 = (((downsize_d_sel ^ 1'b0) & _zz_when_WidthAdapter_l84) == 1'b0);
  assign when_WidthAdapter_l84_1 = (((downsize_d_sel ^ 1'b1) & _zz_when_WidthAdapter_l84) == 1'b0);
  always @(posedge litex_clk or posedge litex_reset) begin
    if(litex_reset) begin
      downsize_a_ctrl_counter <= 1'b0;
      io_down_a_tracker_beat <= 4'b0000;
      io_down_d_tracker_beat <= 4'b0000;
      downsize_d_ctrl_buffer_valid <= 1'b0;
      downsize_d_ctrl_buffer_first <= 1'b1;
    end else begin
      if(io_down_a_fire) begin
        io_down_a_tracker_beat <= (io_down_a_tracker_beat + 4'b0001);
        if(downsize_a_ctrl_burstLast) begin
          io_down_a_tracker_beat <= 4'b0000;
        end
      end
      if(io_down_a_fire) begin
        downsize_a_ctrl_counter <= (downsize_a_ctrl_counter + 1'b1);
        if(downsize_a_ctrl_burstLast) begin
          downsize_a_ctrl_counter <= 1'b0;
        end
      end
      if(io_down_d_fire) begin
        io_down_d_tracker_beat <= (io_down_d_tracker_beat + 4'b0001);
        if(downsize_d_ctrl_burstLast) begin
          io_down_d_tracker_beat <= 4'b0000;
        end
      end
      if(io_up_d_ready) begin
        downsize_d_ctrl_buffer_valid <= 1'b0;
      end
      if(io_down_d_fire) begin
        downsize_d_ctrl_buffer_valid <= downsize_d_ctrl_wordLast;
        downsize_d_ctrl_buffer_first <= downsize_d_ctrl_wordLast;
      end
    end
  end

  always @(posedge litex_clk) begin
    if(io_down_d_fire) begin
      if(downsize_d_ctrl_buffer_first) begin
        downsize_d_ctrl_buffer_args_opcode <= io_down_d_payload_opcode;
        downsize_d_ctrl_buffer_args_param <= io_down_d_payload_param;
        downsize_d_ctrl_buffer_args_source <= io_down_d_payload_source;
        downsize_d_ctrl_buffer_args_size <= io_down_d_payload_size;
        downsize_d_ctrl_buffer_corrupt <= 1'b0;
        downsize_d_ctrl_buffer_denied <= 1'b0;
      end
      if(when_WidthAdapter_l84) begin
        downsize_d_ctrl_buffer_data_0 <= io_down_d_payload_data;
      end
      if(when_WidthAdapter_l84_1) begin
        downsize_d_ctrl_buffer_data_1 <= io_down_d_payload_data;
      end
      if(io_down_d_payload_corrupt) begin
        downsize_d_ctrl_buffer_corrupt <= 1'b1;
      end
      if(io_down_d_payload_denied) begin
        downsize_d_ctrl_buffer_denied <= 1'b1;
      end
    end
  end


endmodule

module WidthAdapter (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [1:0]    io_up_a_payload_source,
  input  wire [31:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [7:0]    io_up_a_payload_mask,
  input  wire [63:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [1:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [63:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_down_a_valid,
  input  wire          io_down_a_ready,
  output wire [2:0]    io_down_a_payload_opcode,
  output wire [2:0]    io_down_a_payload_param,
  output wire [1:0]    io_down_a_payload_source,
  output wire [31:0]   io_down_a_payload_address,
  output wire [2:0]    io_down_a_payload_size,
  output wire [15:0]   io_down_a_payload_mask,
  output wire [127:0]  io_down_a_payload_data,
  output wire          io_down_a_payload_corrupt,
  input  wire          io_down_d_valid,
  output wire          io_down_d_ready,
  input  wire [2:0]    io_down_d_payload_opcode,
  input  wire [2:0]    io_down_d_payload_param,
  input  wire [1:0]    io_down_d_payload_source,
  input  wire [2:0]    io_down_d_payload_size,
  input  wire          io_down_d_payload_denied,
  input  wire [127:0]  io_down_d_payload_data,
  input  wire          io_down_d_payload_corrupt,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                upsize_d_ctx_io_add_valid;
  wire       [0:0]    upsize_d_ctx_io_add_payload_context;
  wire                upsize_d_ctx_io_remove_valid;
  wire                upsize_d_ctx_io_add_ready;
  wire       [0:0]    upsize_d_ctx_io_query_context;
  reg        [2:0]    _zz_upsize_a_ctrl_burstLast;
  reg        [2:0]    _zz_io_up_a_tracker_last;
  reg        [2:0]    _zz_upsize_d_ctrl_burstLast;
  reg        [63:0]   _zz_io_up_d_payload_data;
  reg                 upsize_iaHalt;
  wire                _zz_io_up_a_ready;
  wire                upsize_ia_valid;
  wire                upsize_ia_ready;
  wire       [2:0]    upsize_ia_payload_opcode;
  wire       [2:0]    upsize_ia_payload_param;
  wire       [1:0]    upsize_ia_payload_source;
  wire       [31:0]   upsize_ia_payload_address;
  wire       [2:0]    upsize_ia_payload_size;
  wire       [7:0]    upsize_ia_payload_mask;
  wire       [63:0]   upsize_ia_payload_data;
  wire                upsize_ia_payload_corrupt;
  wire       [0:0]    _zz_upsize_a_ctrl_wordLast;
  reg        [2:0]    upsize_ia_tracker_beat;
  wire                upsize_a_ctrl_burstLast;
  wire                upsize_ia_fire;
  wire                upsize_a_ctrl_wordLast;
  reg                 upsize_a_ctrl_buffer_valid;
  reg                 upsize_a_ctrl_buffer_first;
  reg        [2:0]    upsize_a_ctrl_buffer_args_opcode;
  reg        [2:0]    upsize_a_ctrl_buffer_args_param;
  reg        [1:0]    upsize_a_ctrl_buffer_args_source;
  reg        [31:0]   upsize_a_ctrl_buffer_args_address;
  reg        [2:0]    upsize_a_ctrl_buffer_args_size;
  reg        [63:0]   upsize_a_ctrl_buffer_data_0;
  reg        [63:0]   upsize_a_ctrl_buffer_data_1;
  reg        [7:0]    upsize_a_ctrl_buffer_mask_0;
  reg        [7:0]    upsize_a_ctrl_buffer_mask_1;
  reg                 upsize_a_ctrl_buffer_corrupt;
  wire       [1:0]    _zz_1;
  wire       [1:0]    _zz_2;
  wire                io_up_a_fire;
  reg        [2:0]    io_up_a_tracker_beat;
  wire                io_up_a_tracker_last;
  wire                when_ContextBuffer_l19;
  wire                io_up_d_fire;
  reg        [2:0]    io_up_d_tracker_beat;
  wire                upsize_d_ctrl_burstLast;
  reg        [0:0]    upsize_d_ctrl_counter;
  wire       [0:0]    upsize_d_ctrl_sel;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] io_down_a_payload_opcode_string;
  reg [119:0] io_down_d_payload_opcode_string;
  reg [127:0] upsize_ia_payload_opcode_string;
  reg [127:0] upsize_a_ctrl_buffer_args_opcode_string;
  `endif


  ContextAsyncBufferFull_1 upsize_d_ctx (
    .io_add_valid           (upsize_d_ctx_io_add_valid          ), //i
    .io_add_ready           (upsize_d_ctx_io_add_ready          ), //o
    .io_add_payload_id      (io_up_a_payload_source[1:0]        ), //i
    .io_add_payload_context (upsize_d_ctx_io_add_payload_context), //i
    .io_remove_valid        (upsize_d_ctx_io_remove_valid       ), //i
    .io_remove_payload_id   (io_up_d_payload_source[1:0]        ), //i
    .io_query_id            (io_down_d_payload_source[1:0]      ), //i
    .io_query_context       (upsize_d_ctx_io_query_context      ), //o
    .litex_clk              (litex_clk                          )  //i
  );
  always @(*) begin
    case(upsize_ia_payload_size)
      3'b000 : _zz_upsize_a_ctrl_burstLast = 3'b000;
      3'b001 : _zz_upsize_a_ctrl_burstLast = 3'b000;
      3'b010 : _zz_upsize_a_ctrl_burstLast = 3'b000;
      3'b011 : _zz_upsize_a_ctrl_burstLast = 3'b000;
      3'b100 : _zz_upsize_a_ctrl_burstLast = 3'b001;
      3'b101 : _zz_upsize_a_ctrl_burstLast = 3'b011;
      default : _zz_upsize_a_ctrl_burstLast = 3'b111;
    endcase
  end

  always @(*) begin
    case(io_up_a_payload_size)
      3'b000 : _zz_io_up_a_tracker_last = 3'b000;
      3'b001 : _zz_io_up_a_tracker_last = 3'b000;
      3'b010 : _zz_io_up_a_tracker_last = 3'b000;
      3'b011 : _zz_io_up_a_tracker_last = 3'b000;
      3'b100 : _zz_io_up_a_tracker_last = 3'b001;
      3'b101 : _zz_io_up_a_tracker_last = 3'b011;
      default : _zz_io_up_a_tracker_last = 3'b111;
    endcase
  end

  always @(*) begin
    case(io_up_d_payload_size)
      3'b000 : _zz_upsize_d_ctrl_burstLast = 3'b000;
      3'b001 : _zz_upsize_d_ctrl_burstLast = 3'b000;
      3'b010 : _zz_upsize_d_ctrl_burstLast = 3'b000;
      3'b011 : _zz_upsize_d_ctrl_burstLast = 3'b000;
      3'b100 : _zz_upsize_d_ctrl_burstLast = 3'b001;
      3'b101 : _zz_upsize_d_ctrl_burstLast = 3'b011;
      default : _zz_upsize_d_ctrl_burstLast = 3'b111;
    endcase
  end

  always @(*) begin
    case(upsize_d_ctrl_sel)
      1'b0 : _zz_io_up_d_payload_data = io_down_d_payload_data[63 : 0];
      default : _zz_io_up_d_payload_data = io_down_d_payload_data[127 : 64];
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_down_a_payload_opcode)
      A_PUT_FULL_DATA : io_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_down_d_payload_opcode)
      D_ACCESS_ACK : io_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(upsize_ia_payload_opcode)
      A_PUT_FULL_DATA : upsize_ia_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : upsize_ia_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : upsize_ia_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : upsize_ia_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : upsize_ia_payload_opcode_string = "ACQUIRE_PERM    ";
      default : upsize_ia_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(upsize_a_ctrl_buffer_args_opcode)
      A_PUT_FULL_DATA : upsize_a_ctrl_buffer_args_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : upsize_a_ctrl_buffer_args_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : upsize_a_ctrl_buffer_args_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : upsize_a_ctrl_buffer_args_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : upsize_a_ctrl_buffer_args_opcode_string = "ACQUIRE_PERM    ";
      default : upsize_a_ctrl_buffer_args_opcode_string = "????????????????";
    endcase
  end
  `endif

  always @(*) begin
    upsize_iaHalt = 1'b0;
    if(when_ContextBuffer_l19) begin
      upsize_iaHalt = 1'b1;
    end
  end

  assign _zz_io_up_a_ready = (! upsize_iaHalt);
  assign upsize_ia_valid = (io_up_a_valid && _zz_io_up_a_ready);
  assign io_up_a_ready = (upsize_ia_ready && _zz_io_up_a_ready);
  assign upsize_ia_payload_opcode = io_up_a_payload_opcode;
  assign upsize_ia_payload_param = io_up_a_payload_param;
  assign upsize_ia_payload_source = io_up_a_payload_source;
  assign upsize_ia_payload_address = io_up_a_payload_address;
  assign upsize_ia_payload_size = io_up_a_payload_size;
  assign upsize_ia_payload_mask = io_up_a_payload_mask;
  assign upsize_ia_payload_data = io_up_a_payload_data;
  assign upsize_ia_payload_corrupt = io_up_a_payload_corrupt;
  assign _zz_upsize_a_ctrl_wordLast = upsize_ia_payload_address[3 : 3];
  assign upsize_a_ctrl_burstLast = ((! ((1'b0 || (A_PUT_FULL_DATA == upsize_ia_payload_opcode)) || (A_PUT_PARTIAL_DATA == upsize_ia_payload_opcode))) || (upsize_ia_tracker_beat == _zz_upsize_a_ctrl_burstLast));
  assign upsize_ia_fire = (upsize_ia_valid && upsize_ia_ready);
  assign upsize_a_ctrl_wordLast = ((&_zz_upsize_a_ctrl_wordLast) || upsize_a_ctrl_burstLast);
  assign io_down_a_valid = upsize_a_ctrl_buffer_valid;
  assign io_down_a_payload_opcode = upsize_a_ctrl_buffer_args_opcode;
  assign io_down_a_payload_param = upsize_a_ctrl_buffer_args_param;
  assign io_down_a_payload_source = upsize_a_ctrl_buffer_args_source;
  assign io_down_a_payload_address = upsize_a_ctrl_buffer_args_address;
  assign io_down_a_payload_size = upsize_a_ctrl_buffer_args_size;
  assign io_down_a_payload_mask = {upsize_a_ctrl_buffer_mask_1,upsize_a_ctrl_buffer_mask_0};
  assign io_down_a_payload_data = {upsize_a_ctrl_buffer_data_1,upsize_a_ctrl_buffer_data_0};
  assign io_down_a_payload_corrupt = upsize_a_ctrl_buffer_corrupt;
  assign upsize_ia_ready = ((! upsize_a_ctrl_buffer_valid) || io_down_a_ready);
  assign _zz_1 = ({1'd0,1'b1} <<< _zz_upsize_a_ctrl_wordLast);
  assign _zz_2 = ({1'd0,1'b1} <<< _zz_upsize_a_ctrl_wordLast);
  assign io_up_a_fire = (io_up_a_valid && io_up_a_ready);
  assign io_up_a_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == io_up_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_up_a_payload_opcode))) || (io_up_a_tracker_beat == _zz_io_up_a_tracker_last));
  assign upsize_d_ctx_io_add_valid = (io_up_a_fire && io_up_a_tracker_last);
  assign when_ContextBuffer_l19 = (! upsize_d_ctx_io_add_ready);
  assign io_up_d_fire = (io_up_d_valid && io_up_d_ready);
  assign upsize_d_ctrl_burstLast = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_up_d_payload_opcode)) || (D_GRANT_DATA == io_up_d_payload_opcode))) || (io_up_d_tracker_beat == _zz_upsize_d_ctrl_burstLast));
  assign upsize_d_ctx_io_remove_valid = ((io_up_d_fire && upsize_d_ctrl_burstLast) && (|{(io_up_d_payload_opcode == D_GRANT_DATA),{(io_up_d_payload_opcode == D_GRANT),{(io_up_d_payload_opcode == D_ACCESS_ACK_DATA),(io_up_d_payload_opcode == D_ACCESS_ACK)}}}));
  assign upsize_d_ctx_io_add_payload_context = io_up_a_payload_address[3 : 3];
  assign upsize_d_ctrl_sel = (upsize_d_ctrl_counter + upsize_d_ctx_io_query_context);
  assign io_up_d_valid = io_down_d_valid;
  assign io_up_d_payload_opcode = io_down_d_payload_opcode;
  assign io_up_d_payload_param = io_down_d_payload_param;
  assign io_up_d_payload_source = io_down_d_payload_source;
  assign io_up_d_payload_size = io_down_d_payload_size;
  assign io_up_d_payload_denied = io_down_d_payload_denied;
  assign io_up_d_payload_corrupt = io_down_d_payload_corrupt;
  assign io_down_d_ready = (io_up_d_ready && ((&upsize_d_ctrl_counter) || upsize_d_ctrl_burstLast));
  assign io_up_d_payload_data = _zz_io_up_d_payload_data;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      upsize_ia_tracker_beat <= 3'b000;
      upsize_a_ctrl_buffer_valid <= 1'b0;
      upsize_a_ctrl_buffer_first <= 1'b1;
      io_up_a_tracker_beat <= 3'b000;
      io_up_d_tracker_beat <= 3'b000;
      upsize_d_ctrl_counter <= 1'b0;
    end else begin
      if(upsize_ia_fire) begin
        upsize_ia_tracker_beat <= (upsize_ia_tracker_beat + 3'b001);
        if(upsize_a_ctrl_burstLast) begin
          upsize_ia_tracker_beat <= 3'b000;
        end
      end
      if(io_down_a_ready) begin
        upsize_a_ctrl_buffer_valid <= 1'b0;
      end
      if(upsize_ia_fire) begin
        upsize_a_ctrl_buffer_valid <= upsize_a_ctrl_wordLast;
        upsize_a_ctrl_buffer_first <= upsize_a_ctrl_wordLast;
      end
      if(io_up_a_fire) begin
        io_up_a_tracker_beat <= (io_up_a_tracker_beat + 3'b001);
        if(io_up_a_tracker_last) begin
          io_up_a_tracker_beat <= 3'b000;
        end
      end
      if(io_up_d_fire) begin
        io_up_d_tracker_beat <= (io_up_d_tracker_beat + 3'b001);
        if(upsize_d_ctrl_burstLast) begin
          io_up_d_tracker_beat <= 3'b000;
        end
      end
      if(io_up_d_fire) begin
        upsize_d_ctrl_counter <= (upsize_d_ctrl_counter + 1'b1);
        if(upsize_d_ctrl_burstLast) begin
          upsize_d_ctrl_counter <= 1'b0;
        end
      end
    end
  end

  always @(posedge litex_clk) begin
    if(upsize_ia_fire) begin
      if(upsize_a_ctrl_buffer_first) begin
        upsize_a_ctrl_buffer_args_opcode <= upsize_ia_payload_opcode;
        upsize_a_ctrl_buffer_args_param <= upsize_ia_payload_param;
        upsize_a_ctrl_buffer_args_source <= upsize_ia_payload_source;
        upsize_a_ctrl_buffer_args_address <= upsize_ia_payload_address;
        upsize_a_ctrl_buffer_args_size <= upsize_ia_payload_size;
        upsize_a_ctrl_buffer_corrupt <= 1'b0;
        upsize_a_ctrl_buffer_mask_0 <= 8'h0;
        upsize_a_ctrl_buffer_mask_1 <= 8'h0;
      end
      if(_zz_1[0]) begin
        upsize_a_ctrl_buffer_data_0 <= upsize_ia_payload_data;
      end
      if(_zz_1[1]) begin
        upsize_a_ctrl_buffer_data_1 <= upsize_ia_payload_data;
      end
      if(_zz_2[0]) begin
        upsize_a_ctrl_buffer_mask_0 <= upsize_ia_payload_mask;
      end
      if(_zz_2[1]) begin
        upsize_a_ctrl_buffer_mask_1 <= upsize_ia_payload_mask;
      end
      if(upsize_ia_payload_corrupt) begin
        upsize_a_ctrl_buffer_corrupt <= 1'b1;
      end
    end
  end


endmodule

module AxiLite4Bridge (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [2:0]    io_up_a_payload_source,
  input  wire [31:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [3:0]    io_up_a_payload_mask,
  input  wire [31:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [2:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [31:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_down_aw_valid,
  input  wire          io_down_aw_ready,
  output wire [31:0]   io_down_aw_payload_addr,
  output wire [2:0]    io_down_aw_payload_prot,
  output wire          io_down_w_valid,
  input  wire          io_down_w_ready,
  output wire [31:0]   io_down_w_payload_data,
  output wire [3:0]    io_down_w_payload_strb,
  input  wire          io_down_b_valid,
  output wire          io_down_b_ready,
  input  wire [1:0]    io_down_b_payload_resp,
  output wire          io_down_ar_valid,
  input  wire          io_down_ar_ready,
  output wire [31:0]   io_down_ar_payload_addr,
  output wire [2:0]    io_down_ar_payload_prot,
  input  wire          io_down_r_valid,
  output wire          io_down_r_ready,
  input  wire [31:0]   io_down_r_payload_data,
  input  wire [1:0]    io_down_r_payload_resp,
  input  wire          litex_clk,
  input  wire          litex_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  reg        [3:0]    _zz__zz_io_up_d_tracker_last;
  reg        [3:0]    _zz_io_up_a_tracker_last;
  reg        [3:0]    _zz_a_cmdFork_ready;
  wire       [31:0]   _zz_a_cmd_address;
  wire       [5:0]    _zz_a_cmd_address_1;
  reg                 pending_valid;
  wire                io_up_d_fire;
  reg        [3:0]    io_up_d_tracker_beat;
  wire       [3:0]    _zz_io_up_d_tracker_last;
  wire                io_up_d_tracker_last;
  wire                when_AxiLite4Bridge_l29;
  reg                 pending_get;
  reg        [2:0]    pending_source;
  reg        [2:0]    pending_size;
  reg        [3:0]    io_up_a_tracker_beat;
  wire                io_up_a_tracker_last;
  wire                io_up_a_fire;
  wire                _zz_io_up_a_ready;
  wire                a_halted_valid;
  wire                a_halted_ready;
  wire       [2:0]    a_halted_payload_opcode;
  wire       [2:0]    a_halted_payload_param;
  wire       [2:0]    a_halted_payload_source;
  wire       [31:0]   a_halted_payload_address;
  wire       [2:0]    a_halted_payload_size;
  wire       [3:0]    a_halted_payload_mask;
  wire       [31:0]   a_halted_payload_data;
  wire                a_halted_payload_corrupt;
  wire                a_halted_fire;
  wire                a_buffered_valid;
  reg                 a_buffered_ready;
  wire       [2:0]    a_buffered_payload_opcode;
  wire       [2:0]    a_buffered_payload_param;
  wire       [2:0]    a_buffered_payload_source;
  wire       [31:0]   a_buffered_payload_address;
  wire       [2:0]    a_buffered_payload_size;
  wire       [3:0]    a_buffered_payload_mask;
  wire       [31:0]   a_buffered_payload_data;
  wire                a_buffered_payload_corrupt;
  reg                 a_halted_rValid;
  wire                a_buffered_fire;
  reg        [2:0]    a_halted_rData_opcode;
  reg        [2:0]    a_halted_rData_param;
  reg        [2:0]    a_halted_rData_source;
  reg        [31:0]   a_halted_rData_address;
  reg        [2:0]    a_halted_rData_size;
  reg        [3:0]    a_halted_rData_mask;
  reg        [31:0]   a_halted_rData_data;
  reg                 a_halted_rData_corrupt;
  wire                a_cmdFork_valid;
  wire                a_cmdFork_ready;
  wire       [2:0]    a_cmdFork_payload_opcode;
  wire       [2:0]    a_cmdFork_payload_param;
  wire       [2:0]    a_cmdFork_payload_source;
  wire       [31:0]   a_cmdFork_payload_address;
  wire       [2:0]    a_cmdFork_payload_size;
  wire       [3:0]    a_cmdFork_payload_mask;
  wire       [31:0]   a_cmdFork_payload_data;
  wire                a_cmdFork_payload_corrupt;
  wire                a_dataFork_valid;
  reg                 a_dataFork_ready;
  wire       [2:0]    a_dataFork_payload_opcode;
  wire       [2:0]    a_dataFork_payload_param;
  wire       [2:0]    a_dataFork_payload_source;
  wire       [31:0]   a_dataFork_payload_address;
  wire       [2:0]    a_dataFork_payload_size;
  wire       [3:0]    a_dataFork_payload_mask;
  wire       [31:0]   a_dataFork_payload_data;
  wire                a_dataFork_payload_corrupt;
  reg                 a_buffered_fork2_logic_linkEnable_0;
  reg                 a_buffered_fork2_logic_linkEnable_1;
  wire                when_Stream_l1094;
  wire                when_Stream_l1094_1;
  wire                a_cmdFork_fire;
  wire                a_dataFork_fire;
  wire                a_cmd_isGet;
  reg        [3:0]    a_cmd_counter;
  wire                a_cmd_forked_valid;
  wire                a_cmd_forked_ready;
  wire       [2:0]    a_cmd_forked_payload_opcode;
  wire       [2:0]    a_cmd_forked_payload_param;
  wire       [2:0]    a_cmd_forked_payload_source;
  wire       [31:0]   a_cmd_forked_payload_address;
  wire       [2:0]    a_cmd_forked_payload_size;
  wire       [3:0]    a_cmd_forked_payload_mask;
  wire       [31:0]   a_cmd_forked_payload_data;
  wire                a_cmd_forked_payload_corrupt;
  wire                a_cmd_forked_fire;
  wire       [31:0]   a_cmd_address;
  wire                when_Stream_l472;
  reg                 a_data_filtred_valid;
  wire                a_data_filtred_ready;
  wire       [2:0]    a_data_filtred_payload_opcode;
  wire       [2:0]    a_data_filtred_payload_param;
  wire       [2:0]    a_data_filtred_payload_source;
  wire       [31:0]   a_data_filtred_payload_address;
  wire       [2:0]    a_data_filtred_payload_size;
  wire       [3:0]    a_data_filtred_payload_mask;
  wire       [31:0]   a_data_filtred_payload_data;
  wire                a_data_filtred_payload_corrupt;
  reg        [3:0]    d_counter;
  wire                d_lastB;
  wire                io_down_b_fire;
  wire       [2:0]    _zz_io_up_d_payload_opcode;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] a_halted_payload_opcode_string;
  reg [127:0] a_buffered_payload_opcode_string;
  reg [127:0] a_halted_rData_opcode_string;
  reg [127:0] a_cmdFork_payload_opcode_string;
  reg [127:0] a_dataFork_payload_opcode_string;
  reg [127:0] a_cmd_forked_payload_opcode_string;
  reg [127:0] a_data_filtred_payload_opcode_string;
  reg [119:0] _zz_io_up_d_payload_opcode_string;
  `endif


  assign _zz_a_cmd_address_1 = ({2'd0,a_cmd_counter} <<< 2'd2);
  assign _zz_a_cmd_address = {26'd0, _zz_a_cmd_address_1};
  always @(*) begin
    case(io_up_d_payload_size)
      3'b000 : _zz__zz_io_up_d_tracker_last = 4'b0000;
      3'b001 : _zz__zz_io_up_d_tracker_last = 4'b0000;
      3'b010 : _zz__zz_io_up_d_tracker_last = 4'b0000;
      3'b011 : _zz__zz_io_up_d_tracker_last = 4'b0001;
      3'b100 : _zz__zz_io_up_d_tracker_last = 4'b0011;
      3'b101 : _zz__zz_io_up_d_tracker_last = 4'b0111;
      default : _zz__zz_io_up_d_tracker_last = 4'b1111;
    endcase
  end

  always @(*) begin
    case(io_up_a_payload_size)
      3'b000 : _zz_io_up_a_tracker_last = 4'b0000;
      3'b001 : _zz_io_up_a_tracker_last = 4'b0000;
      3'b010 : _zz_io_up_a_tracker_last = 4'b0000;
      3'b011 : _zz_io_up_a_tracker_last = 4'b0001;
      3'b100 : _zz_io_up_a_tracker_last = 4'b0011;
      3'b101 : _zz_io_up_a_tracker_last = 4'b0111;
      default : _zz_io_up_a_tracker_last = 4'b1111;
    endcase
  end

  always @(*) begin
    case(a_cmdFork_payload_size)
      3'b000 : _zz_a_cmdFork_ready = 4'b0000;
      3'b001 : _zz_a_cmdFork_ready = 4'b0000;
      3'b010 : _zz_a_cmdFork_ready = 4'b0000;
      3'b011 : _zz_a_cmdFork_ready = 4'b0001;
      3'b100 : _zz_a_cmdFork_ready = 4'b0011;
      3'b101 : _zz_a_cmdFork_ready = 4'b0111;
      default : _zz_a_cmdFork_ready = 4'b1111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(a_halted_payload_opcode)
      A_PUT_FULL_DATA : a_halted_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_halted_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_halted_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_halted_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_halted_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_halted_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_buffered_payload_opcode)
      A_PUT_FULL_DATA : a_buffered_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_buffered_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_buffered_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_buffered_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_buffered_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_buffered_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_halted_rData_opcode)
      A_PUT_FULL_DATA : a_halted_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_halted_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_halted_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_halted_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_halted_rData_opcode_string = "ACQUIRE_PERM    ";
      default : a_halted_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmdFork_payload_opcode)
      A_PUT_FULL_DATA : a_cmdFork_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmdFork_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmdFork_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmdFork_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmdFork_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmdFork_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_dataFork_payload_opcode)
      A_PUT_FULL_DATA : a_dataFork_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_dataFork_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_dataFork_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_dataFork_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_dataFork_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_dataFork_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmd_forked_payload_opcode)
      A_PUT_FULL_DATA : a_cmd_forked_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmd_forked_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmd_forked_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmd_forked_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmd_forked_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmd_forked_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_data_filtred_payload_opcode)
      A_PUT_FULL_DATA : a_data_filtred_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_data_filtred_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_data_filtred_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_data_filtred_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_data_filtred_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_data_filtred_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_d_payload_opcode)
      D_ACCESS_ACK : _zz_io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign io_up_d_fire = (io_up_d_valid && io_up_d_ready);
  assign _zz_io_up_d_tracker_last = _zz__zz_io_up_d_tracker_last;
  assign io_up_d_tracker_last = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_up_d_payload_opcode)) || (D_GRANT_DATA == io_up_d_payload_opcode))) || (io_up_d_tracker_beat == _zz_io_up_d_tracker_last));
  assign when_AxiLite4Bridge_l29 = (io_up_d_fire && io_up_d_tracker_last);
  assign io_up_a_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == io_up_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_up_a_payload_opcode))) || (io_up_a_tracker_beat == _zz_io_up_a_tracker_last));
  assign io_up_a_fire = (io_up_a_valid && io_up_a_ready);
  assign _zz_io_up_a_ready = (! (pending_valid && (io_up_a_tracker_beat == 4'b0000)));
  assign a_halted_valid = (io_up_a_valid && _zz_io_up_a_ready);
  assign io_up_a_ready = (a_halted_ready && _zz_io_up_a_ready);
  assign a_halted_payload_opcode = io_up_a_payload_opcode;
  assign a_halted_payload_param = io_up_a_payload_param;
  assign a_halted_payload_source = io_up_a_payload_source;
  assign a_halted_payload_address = io_up_a_payload_address;
  assign a_halted_payload_size = io_up_a_payload_size;
  assign a_halted_payload_mask = io_up_a_payload_mask;
  assign a_halted_payload_data = io_up_a_payload_data;
  assign a_halted_payload_corrupt = io_up_a_payload_corrupt;
  assign a_halted_fire = (a_halted_valid && a_halted_ready);
  assign a_buffered_fire = (a_buffered_valid && a_buffered_ready);
  assign a_halted_ready = (! a_halted_rValid);
  assign a_buffered_valid = a_halted_rValid;
  assign a_buffered_payload_opcode = a_halted_rData_opcode;
  assign a_buffered_payload_param = a_halted_rData_param;
  assign a_buffered_payload_source = a_halted_rData_source;
  assign a_buffered_payload_address = a_halted_rData_address;
  assign a_buffered_payload_size = a_halted_rData_size;
  assign a_buffered_payload_mask = a_halted_rData_mask;
  assign a_buffered_payload_data = a_halted_rData_data;
  assign a_buffered_payload_corrupt = a_halted_rData_corrupt;
  always @(*) begin
    a_buffered_ready = 1'b1;
    if(when_Stream_l1094) begin
      a_buffered_ready = 1'b0;
    end
    if(when_Stream_l1094_1) begin
      a_buffered_ready = 1'b0;
    end
  end

  assign when_Stream_l1094 = ((! a_cmdFork_ready) && a_buffered_fork2_logic_linkEnable_0);
  assign when_Stream_l1094_1 = ((! a_dataFork_ready) && a_buffered_fork2_logic_linkEnable_1);
  assign a_cmdFork_valid = (a_buffered_valid && a_buffered_fork2_logic_linkEnable_0);
  assign a_cmdFork_payload_opcode = a_buffered_payload_opcode;
  assign a_cmdFork_payload_param = a_buffered_payload_param;
  assign a_cmdFork_payload_source = a_buffered_payload_source;
  assign a_cmdFork_payload_address = a_buffered_payload_address;
  assign a_cmdFork_payload_size = a_buffered_payload_size;
  assign a_cmdFork_payload_mask = a_buffered_payload_mask;
  assign a_cmdFork_payload_data = a_buffered_payload_data;
  assign a_cmdFork_payload_corrupt = a_buffered_payload_corrupt;
  assign a_cmdFork_fire = (a_cmdFork_valid && a_cmdFork_ready);
  assign a_dataFork_valid = (a_buffered_valid && a_buffered_fork2_logic_linkEnable_1);
  assign a_dataFork_payload_opcode = a_buffered_payload_opcode;
  assign a_dataFork_payload_param = a_buffered_payload_param;
  assign a_dataFork_payload_source = a_buffered_payload_source;
  assign a_dataFork_payload_address = a_buffered_payload_address;
  assign a_dataFork_payload_size = a_buffered_payload_size;
  assign a_dataFork_payload_mask = a_buffered_payload_mask;
  assign a_dataFork_payload_data = a_buffered_payload_data;
  assign a_dataFork_payload_corrupt = a_buffered_payload_corrupt;
  assign a_dataFork_fire = (a_dataFork_valid && a_dataFork_ready);
  assign a_cmd_isGet = (a_cmdFork_payload_opcode == A_GET);
  assign a_cmd_forked_valid = a_cmdFork_valid;
  assign a_cmd_forked_payload_opcode = a_cmdFork_payload_opcode;
  assign a_cmd_forked_payload_param = a_cmdFork_payload_param;
  assign a_cmd_forked_payload_source = a_cmdFork_payload_source;
  assign a_cmd_forked_payload_address = a_cmdFork_payload_address;
  assign a_cmd_forked_payload_size = a_cmdFork_payload_size;
  assign a_cmd_forked_payload_mask = a_cmdFork_payload_mask;
  assign a_cmd_forked_payload_data = a_cmdFork_payload_data;
  assign a_cmd_forked_payload_corrupt = a_cmdFork_payload_corrupt;
  assign a_cmdFork_ready = (a_cmd_forked_ready && ((! a_cmd_isGet) || (a_cmd_counter == _zz_a_cmdFork_ready)));
  assign a_cmd_forked_fire = (a_cmd_forked_valid && a_cmd_forked_ready);
  assign io_down_aw_valid = (a_cmd_forked_valid && (! a_cmd_isGet));
  assign io_down_ar_valid = (a_cmd_forked_valid && a_cmd_isGet);
  assign a_cmd_forked_ready = (a_cmd_isGet ? io_down_ar_ready : io_down_aw_ready);
  assign a_cmd_address = (a_cmd_forked_payload_address | _zz_a_cmd_address);
  assign io_down_aw_payload_addr = a_cmd_address;
  assign io_down_aw_payload_prot = 3'b010;
  assign io_down_ar_payload_addr = a_cmd_address;
  assign io_down_ar_payload_prot = 3'b010;
  assign when_Stream_l472 = (! ((a_dataFork_payload_opcode == A_PUT_FULL_DATA) || (a_dataFork_payload_opcode == A_PUT_PARTIAL_DATA)));
  always @(*) begin
    a_data_filtred_valid = a_dataFork_valid;
    if(when_Stream_l472) begin
      a_data_filtred_valid = 1'b0;
    end
  end

  always @(*) begin
    a_dataFork_ready = a_data_filtred_ready;
    if(when_Stream_l472) begin
      a_dataFork_ready = 1'b1;
    end
  end

  assign a_data_filtred_payload_opcode = a_dataFork_payload_opcode;
  assign a_data_filtred_payload_param = a_dataFork_payload_param;
  assign a_data_filtred_payload_source = a_dataFork_payload_source;
  assign a_data_filtred_payload_address = a_dataFork_payload_address;
  assign a_data_filtred_payload_size = a_dataFork_payload_size;
  assign a_data_filtred_payload_mask = a_dataFork_payload_mask;
  assign a_data_filtred_payload_data = a_dataFork_payload_data;
  assign a_data_filtred_payload_corrupt = a_dataFork_payload_corrupt;
  assign io_down_w_valid = a_data_filtred_valid;
  assign a_data_filtred_ready = io_down_w_ready;
  assign io_down_w_payload_data = a_data_filtred_payload_data;
  assign io_down_w_payload_strb = a_data_filtred_payload_mask;
  assign d_lastB = (d_counter == _zz_io_up_d_tracker_last);
  assign io_down_b_fire = (io_down_b_valid && io_down_b_ready);
  assign io_down_r_ready = io_up_d_ready;
  assign io_down_b_ready = (io_up_d_ready || (! d_lastB));
  assign io_up_d_valid = (io_down_r_valid || (io_down_b_valid && d_lastB));
  assign _zz_io_up_d_payload_opcode = (pending_get ? D_ACCESS_ACK_DATA : D_ACCESS_ACK);
  assign io_up_d_payload_opcode = _zz_io_up_d_payload_opcode;
  assign io_up_d_payload_param = 3'b000;
  assign io_up_d_payload_source = pending_source;
  assign io_up_d_payload_denied = (! (pending_get ? (io_down_r_payload_resp == 2'b00) : (io_down_b_payload_resp == 2'b00)));
  assign io_up_d_payload_data = io_down_r_payload_data;
  assign io_up_d_payload_corrupt = 1'b0;
  assign io_up_d_payload_size = pending_size;
  always @(posedge litex_clk or posedge litex_reset) begin
    if(litex_reset) begin
      pending_valid <= 1'b0;
      io_up_d_tracker_beat <= 4'b0000;
      io_up_a_tracker_beat <= 4'b0000;
      a_halted_rValid <= 1'b0;
      a_buffered_fork2_logic_linkEnable_0 <= 1'b1;
      a_buffered_fork2_logic_linkEnable_1 <= 1'b1;
      a_cmd_counter <= 4'b0000;
      d_counter <= 4'b0000;
    end else begin
      if(io_up_d_fire) begin
        io_up_d_tracker_beat <= (io_up_d_tracker_beat + 4'b0001);
        if(io_up_d_tracker_last) begin
          io_up_d_tracker_beat <= 4'b0000;
        end
      end
      if(when_AxiLite4Bridge_l29) begin
        pending_valid <= 1'b0;
      end
      if(io_up_a_fire) begin
        io_up_a_tracker_beat <= (io_up_a_tracker_beat + 4'b0001);
        if(io_up_a_tracker_last) begin
          io_up_a_tracker_beat <= 4'b0000;
        end
      end
      if(a_halted_fire) begin
        pending_valid <= 1'b1;
      end
      if(a_halted_valid) begin
        a_halted_rValid <= 1'b1;
      end
      if(a_buffered_fire) begin
        a_halted_rValid <= 1'b0;
      end
      if(a_cmdFork_fire) begin
        a_buffered_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(a_dataFork_fire) begin
        a_buffered_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(a_buffered_ready) begin
        a_buffered_fork2_logic_linkEnable_0 <= 1'b1;
        a_buffered_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(a_cmd_forked_fire) begin
        a_cmd_counter <= (a_cmd_counter + 4'b0001);
        if(a_cmdFork_fire) begin
          a_cmd_counter <= 4'b0000;
        end
      end
      if(io_down_b_fire) begin
        d_counter <= (d_counter + 4'b0001);
        if(d_lastB) begin
          d_counter <= 4'b0000;
        end
      end
    end
  end

  always @(posedge litex_clk) begin
    if(a_halted_fire) begin
      pending_get <= (a_halted_payload_opcode == A_GET);
      pending_source <= a_halted_payload_source;
      pending_size <= a_halted_payload_size;
    end
    if(a_halted_ready) begin
      a_halted_rData_opcode <= a_halted_payload_opcode;
      a_halted_rData_param <= a_halted_payload_param;
      a_halted_rData_source <= a_halted_payload_source;
      a_halted_rData_address <= a_halted_payload_address;
      a_halted_rData_size <= a_halted_payload_size;
      a_halted_rData_mask <= a_halted_payload_mask;
      a_halted_rData_data <= a_halted_payload_data;
      a_halted_rData_corrupt <= a_halted_payload_corrupt;
    end
  end


endmodule

module TilelinkPlic (
  input  wire          io_bus_a_valid,
  output wire          io_bus_a_ready,
  input  wire [2:0]    io_bus_a_payload_opcode,
  input  wire [2:0]    io_bus_a_payload_param,
  input  wire [2:0]    io_bus_a_payload_source,
  input  wire [21:0]   io_bus_a_payload_address,
  input  wire [1:0]    io_bus_a_payload_size,
  input  wire [3:0]    io_bus_a_payload_mask,
  input  wire [31:0]   io_bus_a_payload_data,
  input  wire          io_bus_a_payload_corrupt,
  output wire          io_bus_d_valid,
  input  wire          io_bus_d_ready,
  output wire [2:0]    io_bus_d_payload_opcode,
  output wire [2:0]    io_bus_d_payload_param,
  output wire [2:0]    io_bus_d_payload_source,
  output wire [1:0]    io_bus_d_payload_size,
  output wire          io_bus_d_payload_denied,
  output wire [31:0]   io_bus_d_payload_data,
  output wire          io_bus_d_payload_corrupt,
  input  wire [30:0]   io_sources,
  output wire [1:0]    io_targets,
  input  wire          litex_clk,
  input  wire          litex_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire       [4:0]    _zz_targets_0_bestRequest_id_82;
  wire       [4:0]    _zz_targets_0_bestRequest_id_83;
  wire       [4:0]    _zz_targets_0_bestRequest_id_84;
  wire       [4:0]    _zz_targets_0_bestRequest_id_85;
  wire       [4:0]    _zz_targets_0_bestRequest_id_86;
  wire       [4:0]    _zz_targets_0_bestRequest_id_87;
  wire       [4:0]    _zz_targets_0_bestRequest_id_88;
  wire       [4:0]    _zz_targets_0_bestRequest_id_89;
  wire       [4:0]    _zz_targets_0_bestRequest_id_90;
  wire       [4:0]    _zz_targets_0_bestRequest_id_91;
  wire       [4:0]    _zz_targets_0_bestRequest_id_92;
  wire       [4:0]    _zz_targets_0_bestRequest_id_93;
  wire       [4:0]    _zz_targets_0_bestRequest_id_94;
  wire       [4:0]    _zz_targets_0_bestRequest_id_95;
  wire       [4:0]    _zz_targets_0_bestRequest_id_96;
  wire       [4:0]    _zz_targets_0_bestRequest_id_97;
  wire       [4:0]    _zz_targets_1_bestRequest_id_82;
  wire       [4:0]    _zz_targets_1_bestRequest_id_83;
  wire       [4:0]    _zz_targets_1_bestRequest_id_84;
  wire       [4:0]    _zz_targets_1_bestRequest_id_85;
  wire       [4:0]    _zz_targets_1_bestRequest_id_86;
  wire       [4:0]    _zz_targets_1_bestRequest_id_87;
  wire       [4:0]    _zz_targets_1_bestRequest_id_88;
  wire       [4:0]    _zz_targets_1_bestRequest_id_89;
  wire       [4:0]    _zz_targets_1_bestRequest_id_90;
  wire       [4:0]    _zz_targets_1_bestRequest_id_91;
  wire       [4:0]    _zz_targets_1_bestRequest_id_92;
  wire       [4:0]    _zz_targets_1_bestRequest_id_93;
  wire       [4:0]    _zz_targets_1_bestRequest_id_94;
  wire       [4:0]    _zz_targets_1_bestRequest_id_95;
  wire       [4:0]    _zz_targets_1_bestRequest_id_96;
  wire       [4:0]    _zz_targets_1_bestRequest_id_97;
  wire       [19:0]   _zz_factory_address;
  wire                _zz_gateways_0_ip;
  wire                _zz_gateways_1_ip;
  wire                _zz_gateways_2_ip;
  wire                _zz_gateways_3_ip;
  wire                _zz_gateways_4_ip;
  wire                _zz_gateways_5_ip;
  wire                _zz_gateways_6_ip;
  wire                _zz_gateways_7_ip;
  wire                _zz_gateways_8_ip;
  wire                _zz_gateways_9_ip;
  wire                _zz_gateways_10_ip;
  wire                _zz_gateways_11_ip;
  wire                _zz_gateways_12_ip;
  wire                _zz_gateways_13_ip;
  wire                _zz_gateways_14_ip;
  wire                _zz_gateways_15_ip;
  wire                _zz_gateways_16_ip;
  wire                _zz_gateways_17_ip;
  wire                _zz_gateways_18_ip;
  wire                _zz_gateways_19_ip;
  wire                _zz_gateways_20_ip;
  wire                _zz_gateways_21_ip;
  wire                _zz_gateways_22_ip;
  wire                _zz_gateways_23_ip;
  wire                _zz_gateways_24_ip;
  wire                _zz_gateways_25_ip;
  wire                _zz_gateways_26_ip;
  wire                _zz_gateways_27_ip;
  wire                _zz_gateways_28_ip;
  wire                _zz_gateways_29_ip;
  wire                _zz_gateways_30_ip;
  wire       [1:0]    gateways_0_priority;
  reg                 gateways_0_ip;
  reg                 gateways_0_waitCompletion;
  wire                when_PlicGateway_l21;
  wire       [1:0]    gateways_1_priority;
  reg                 gateways_1_ip;
  reg                 gateways_1_waitCompletion;
  wire                when_PlicGateway_l21_1;
  wire       [1:0]    gateways_2_priority;
  reg                 gateways_2_ip;
  reg                 gateways_2_waitCompletion;
  wire                when_PlicGateway_l21_2;
  wire       [1:0]    gateways_3_priority;
  reg                 gateways_3_ip;
  reg                 gateways_3_waitCompletion;
  wire                when_PlicGateway_l21_3;
  wire       [1:0]    gateways_4_priority;
  reg                 gateways_4_ip;
  reg                 gateways_4_waitCompletion;
  wire                when_PlicGateway_l21_4;
  wire       [1:0]    gateways_5_priority;
  reg                 gateways_5_ip;
  reg                 gateways_5_waitCompletion;
  wire                when_PlicGateway_l21_5;
  wire       [1:0]    gateways_6_priority;
  reg                 gateways_6_ip;
  reg                 gateways_6_waitCompletion;
  wire                when_PlicGateway_l21_6;
  wire       [1:0]    gateways_7_priority;
  reg                 gateways_7_ip;
  reg                 gateways_7_waitCompletion;
  wire                when_PlicGateway_l21_7;
  wire       [1:0]    gateways_8_priority;
  reg                 gateways_8_ip;
  reg                 gateways_8_waitCompletion;
  wire                when_PlicGateway_l21_8;
  wire       [1:0]    gateways_9_priority;
  reg                 gateways_9_ip;
  reg                 gateways_9_waitCompletion;
  wire                when_PlicGateway_l21_9;
  wire       [1:0]    gateways_10_priority;
  reg                 gateways_10_ip;
  reg                 gateways_10_waitCompletion;
  wire                when_PlicGateway_l21_10;
  wire       [1:0]    gateways_11_priority;
  reg                 gateways_11_ip;
  reg                 gateways_11_waitCompletion;
  wire                when_PlicGateway_l21_11;
  wire       [1:0]    gateways_12_priority;
  reg                 gateways_12_ip;
  reg                 gateways_12_waitCompletion;
  wire                when_PlicGateway_l21_12;
  wire       [1:0]    gateways_13_priority;
  reg                 gateways_13_ip;
  reg                 gateways_13_waitCompletion;
  wire                when_PlicGateway_l21_13;
  wire       [1:0]    gateways_14_priority;
  reg                 gateways_14_ip;
  reg                 gateways_14_waitCompletion;
  wire                when_PlicGateway_l21_14;
  wire       [1:0]    gateways_15_priority;
  reg                 gateways_15_ip;
  reg                 gateways_15_waitCompletion;
  wire                when_PlicGateway_l21_15;
  wire       [1:0]    gateways_16_priority;
  reg                 gateways_16_ip;
  reg                 gateways_16_waitCompletion;
  wire                when_PlicGateway_l21_16;
  wire       [1:0]    gateways_17_priority;
  reg                 gateways_17_ip;
  reg                 gateways_17_waitCompletion;
  wire                when_PlicGateway_l21_17;
  wire       [1:0]    gateways_18_priority;
  reg                 gateways_18_ip;
  reg                 gateways_18_waitCompletion;
  wire                when_PlicGateway_l21_18;
  wire       [1:0]    gateways_19_priority;
  reg                 gateways_19_ip;
  reg                 gateways_19_waitCompletion;
  wire                when_PlicGateway_l21_19;
  wire       [1:0]    gateways_20_priority;
  reg                 gateways_20_ip;
  reg                 gateways_20_waitCompletion;
  wire                when_PlicGateway_l21_20;
  wire       [1:0]    gateways_21_priority;
  reg                 gateways_21_ip;
  reg                 gateways_21_waitCompletion;
  wire                when_PlicGateway_l21_21;
  wire       [1:0]    gateways_22_priority;
  reg                 gateways_22_ip;
  reg                 gateways_22_waitCompletion;
  wire                when_PlicGateway_l21_22;
  wire       [1:0]    gateways_23_priority;
  reg                 gateways_23_ip;
  reg                 gateways_23_waitCompletion;
  wire                when_PlicGateway_l21_23;
  wire       [1:0]    gateways_24_priority;
  reg                 gateways_24_ip;
  reg                 gateways_24_waitCompletion;
  wire                when_PlicGateway_l21_24;
  wire       [1:0]    gateways_25_priority;
  reg                 gateways_25_ip;
  reg                 gateways_25_waitCompletion;
  wire                when_PlicGateway_l21_25;
  wire       [1:0]    gateways_26_priority;
  reg                 gateways_26_ip;
  reg                 gateways_26_waitCompletion;
  wire                when_PlicGateway_l21_26;
  wire       [1:0]    gateways_27_priority;
  reg                 gateways_27_ip;
  reg                 gateways_27_waitCompletion;
  wire                when_PlicGateway_l21_27;
  wire       [1:0]    gateways_28_priority;
  reg                 gateways_28_ip;
  reg                 gateways_28_waitCompletion;
  wire                when_PlicGateway_l21_28;
  wire       [1:0]    gateways_29_priority;
  reg                 gateways_29_ip;
  reg                 gateways_29_waitCompletion;
  wire                when_PlicGateway_l21_29;
  wire       [1:0]    gateways_30_priority;
  reg                 gateways_30_ip;
  reg                 gateways_30_waitCompletion;
  wire                when_PlicGateway_l21_30;
  wire                targets_0_ie_0;
  wire                targets_0_ie_1;
  wire                targets_0_ie_2;
  wire                targets_0_ie_3;
  wire                targets_0_ie_4;
  wire                targets_0_ie_5;
  wire                targets_0_ie_6;
  wire                targets_0_ie_7;
  wire                targets_0_ie_8;
  wire                targets_0_ie_9;
  wire                targets_0_ie_10;
  wire                targets_0_ie_11;
  wire                targets_0_ie_12;
  wire                targets_0_ie_13;
  wire                targets_0_ie_14;
  wire                targets_0_ie_15;
  wire                targets_0_ie_16;
  wire                targets_0_ie_17;
  wire                targets_0_ie_18;
  wire                targets_0_ie_19;
  wire                targets_0_ie_20;
  wire                targets_0_ie_21;
  wire                targets_0_ie_22;
  wire                targets_0_ie_23;
  wire                targets_0_ie_24;
  wire                targets_0_ie_25;
  wire                targets_0_ie_26;
  wire                targets_0_ie_27;
  wire                targets_0_ie_28;
  wire                targets_0_ie_29;
  wire                targets_0_ie_30;
  wire       [1:0]    targets_0_threshold;
  wire       [1:0]    targets_0_requests_0_priority;
  wire       [4:0]    targets_0_requests_0_id;
  wire                targets_0_requests_0_valid;
  wire       [1:0]    targets_0_requests_1_priority;
  wire       [4:0]    targets_0_requests_1_id;
  wire                targets_0_requests_1_valid;
  wire       [1:0]    targets_0_requests_2_priority;
  wire       [4:0]    targets_0_requests_2_id;
  wire                targets_0_requests_2_valid;
  wire       [1:0]    targets_0_requests_3_priority;
  wire       [4:0]    targets_0_requests_3_id;
  wire                targets_0_requests_3_valid;
  wire       [1:0]    targets_0_requests_4_priority;
  wire       [4:0]    targets_0_requests_4_id;
  wire                targets_0_requests_4_valid;
  wire       [1:0]    targets_0_requests_5_priority;
  wire       [4:0]    targets_0_requests_5_id;
  wire                targets_0_requests_5_valid;
  wire       [1:0]    targets_0_requests_6_priority;
  wire       [4:0]    targets_0_requests_6_id;
  wire                targets_0_requests_6_valid;
  wire       [1:0]    targets_0_requests_7_priority;
  wire       [4:0]    targets_0_requests_7_id;
  wire                targets_0_requests_7_valid;
  wire       [1:0]    targets_0_requests_8_priority;
  wire       [4:0]    targets_0_requests_8_id;
  wire                targets_0_requests_8_valid;
  wire       [1:0]    targets_0_requests_9_priority;
  wire       [4:0]    targets_0_requests_9_id;
  wire                targets_0_requests_9_valid;
  wire       [1:0]    targets_0_requests_10_priority;
  wire       [4:0]    targets_0_requests_10_id;
  wire                targets_0_requests_10_valid;
  wire       [1:0]    targets_0_requests_11_priority;
  wire       [4:0]    targets_0_requests_11_id;
  wire                targets_0_requests_11_valid;
  wire       [1:0]    targets_0_requests_12_priority;
  wire       [4:0]    targets_0_requests_12_id;
  wire                targets_0_requests_12_valid;
  wire       [1:0]    targets_0_requests_13_priority;
  wire       [4:0]    targets_0_requests_13_id;
  wire                targets_0_requests_13_valid;
  wire       [1:0]    targets_0_requests_14_priority;
  wire       [4:0]    targets_0_requests_14_id;
  wire                targets_0_requests_14_valid;
  wire       [1:0]    targets_0_requests_15_priority;
  wire       [4:0]    targets_0_requests_15_id;
  wire                targets_0_requests_15_valid;
  wire       [1:0]    targets_0_requests_16_priority;
  wire       [4:0]    targets_0_requests_16_id;
  wire                targets_0_requests_16_valid;
  wire       [1:0]    targets_0_requests_17_priority;
  wire       [4:0]    targets_0_requests_17_id;
  wire                targets_0_requests_17_valid;
  wire       [1:0]    targets_0_requests_18_priority;
  wire       [4:0]    targets_0_requests_18_id;
  wire                targets_0_requests_18_valid;
  wire       [1:0]    targets_0_requests_19_priority;
  wire       [4:0]    targets_0_requests_19_id;
  wire                targets_0_requests_19_valid;
  wire       [1:0]    targets_0_requests_20_priority;
  wire       [4:0]    targets_0_requests_20_id;
  wire                targets_0_requests_20_valid;
  wire       [1:0]    targets_0_requests_21_priority;
  wire       [4:0]    targets_0_requests_21_id;
  wire                targets_0_requests_21_valid;
  wire       [1:0]    targets_0_requests_22_priority;
  wire       [4:0]    targets_0_requests_22_id;
  wire                targets_0_requests_22_valid;
  wire       [1:0]    targets_0_requests_23_priority;
  wire       [4:0]    targets_0_requests_23_id;
  wire                targets_0_requests_23_valid;
  wire       [1:0]    targets_0_requests_24_priority;
  wire       [4:0]    targets_0_requests_24_id;
  wire                targets_0_requests_24_valid;
  wire       [1:0]    targets_0_requests_25_priority;
  wire       [4:0]    targets_0_requests_25_id;
  wire                targets_0_requests_25_valid;
  wire       [1:0]    targets_0_requests_26_priority;
  wire       [4:0]    targets_0_requests_26_id;
  wire                targets_0_requests_26_valid;
  wire       [1:0]    targets_0_requests_27_priority;
  wire       [4:0]    targets_0_requests_27_id;
  wire                targets_0_requests_27_valid;
  wire       [1:0]    targets_0_requests_28_priority;
  wire       [4:0]    targets_0_requests_28_id;
  wire                targets_0_requests_28_valid;
  wire       [1:0]    targets_0_requests_29_priority;
  wire       [4:0]    targets_0_requests_29_id;
  wire                targets_0_requests_29_valid;
  wire       [1:0]    targets_0_requests_30_priority;
  wire       [4:0]    targets_0_requests_30_id;
  wire                targets_0_requests_30_valid;
  wire       [1:0]    targets_0_requests_31_priority;
  wire       [4:0]    targets_0_requests_31_id;
  wire                targets_0_requests_31_valid;
  wire                _zz_targets_0_bestRequest_id;
  wire       [1:0]    _zz_targets_0_bestRequest_id_1;
  wire                _zz_targets_0_bestRequest_id_2;
  wire                _zz_targets_0_bestRequest_id_3;
  wire       [1:0]    _zz_targets_0_bestRequest_id_4;
  wire                _zz_targets_0_bestRequest_id_5;
  wire                _zz_targets_0_bestRequest_id_6;
  wire       [1:0]    _zz_targets_0_bestRequest_id_7;
  wire                _zz_targets_0_bestRequest_id_8;
  wire                _zz_targets_0_bestRequest_id_9;
  wire       [1:0]    _zz_targets_0_bestRequest_id_10;
  wire                _zz_targets_0_bestRequest_id_11;
  wire                _zz_targets_0_bestRequest_id_12;
  wire       [1:0]    _zz_targets_0_bestRequest_id_13;
  wire                _zz_targets_0_bestRequest_id_14;
  wire                _zz_targets_0_bestRequest_id_15;
  wire       [1:0]    _zz_targets_0_bestRequest_id_16;
  wire                _zz_targets_0_bestRequest_id_17;
  wire                _zz_targets_0_bestRequest_id_18;
  wire       [1:0]    _zz_targets_0_bestRequest_id_19;
  wire                _zz_targets_0_bestRequest_id_20;
  wire                _zz_targets_0_bestRequest_id_21;
  wire       [1:0]    _zz_targets_0_bestRequest_id_22;
  wire                _zz_targets_0_bestRequest_id_23;
  wire                _zz_targets_0_bestRequest_id_24;
  wire       [1:0]    _zz_targets_0_bestRequest_id_25;
  wire                _zz_targets_0_bestRequest_id_26;
  wire                _zz_targets_0_bestRequest_id_27;
  wire       [1:0]    _zz_targets_0_bestRequest_id_28;
  wire                _zz_targets_0_bestRequest_id_29;
  wire                _zz_targets_0_bestRequest_id_30;
  wire       [1:0]    _zz_targets_0_bestRequest_id_31;
  wire                _zz_targets_0_bestRequest_id_32;
  wire                _zz_targets_0_bestRequest_id_33;
  wire       [1:0]    _zz_targets_0_bestRequest_id_34;
  wire                _zz_targets_0_bestRequest_id_35;
  wire                _zz_targets_0_bestRequest_id_36;
  wire       [1:0]    _zz_targets_0_bestRequest_id_37;
  wire                _zz_targets_0_bestRequest_id_38;
  wire                _zz_targets_0_bestRequest_id_39;
  wire       [1:0]    _zz_targets_0_bestRequest_id_40;
  wire                _zz_targets_0_bestRequest_id_41;
  wire                _zz_targets_0_bestRequest_id_42;
  wire       [1:0]    _zz_targets_0_bestRequest_id_43;
  wire                _zz_targets_0_bestRequest_id_44;
  wire                _zz_targets_0_bestRequest_id_45;
  wire       [1:0]    _zz_targets_0_bestRequest_id_46;
  wire                _zz_targets_0_bestRequest_id_47;
  wire                _zz_targets_0_bestRequest_id_48;
  wire       [1:0]    _zz_targets_0_bestRequest_id_49;
  wire                _zz_targets_0_bestRequest_id_50;
  wire                _zz_targets_0_bestRequest_id_51;
  wire       [1:0]    _zz_targets_0_bestRequest_id_52;
  wire                _zz_targets_0_bestRequest_id_53;
  wire                _zz_targets_0_bestRequest_id_54;
  wire       [1:0]    _zz_targets_0_bestRequest_id_55;
  wire                _zz_targets_0_bestRequest_id_56;
  wire                _zz_targets_0_bestRequest_id_57;
  wire       [1:0]    _zz_targets_0_bestRequest_id_58;
  wire                _zz_targets_0_bestRequest_id_59;
  wire                _zz_targets_0_bestRequest_id_60;
  wire       [1:0]    _zz_targets_0_bestRequest_id_61;
  wire                _zz_targets_0_bestRequest_id_62;
  wire                _zz_targets_0_bestRequest_id_63;
  wire       [1:0]    _zz_targets_0_bestRequest_id_64;
  wire                _zz_targets_0_bestRequest_id_65;
  wire                _zz_targets_0_bestRequest_id_66;
  wire       [1:0]    _zz_targets_0_bestRequest_id_67;
  wire                _zz_targets_0_bestRequest_id_68;
  wire                _zz_targets_0_bestRequest_id_69;
  wire       [1:0]    _zz_targets_0_bestRequest_id_70;
  wire                _zz_targets_0_bestRequest_id_71;
  wire                _zz_targets_0_bestRequest_id_72;
  wire       [1:0]    _zz_targets_0_bestRequest_priority;
  wire                _zz_targets_0_bestRequest_id_73;
  wire                _zz_targets_0_bestRequest_id_74;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_1;
  wire                _zz_targets_0_bestRequest_id_75;
  wire                _zz_targets_0_bestRequest_id_76;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_2;
  wire                _zz_targets_0_bestRequest_id_77;
  wire                _zz_targets_0_bestRequest_id_78;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_3;
  wire                _zz_targets_0_bestRequest_id_79;
  wire                _zz_targets_0_bestRequest_id_80;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_4;
  wire                _zz_targets_0_bestRequest_valid;
  wire                _zz_targets_0_bestRequest_id_81;
  wire       [1:0]    _zz_targets_0_bestRequest_priority_5;
  wire                _zz_targets_0_bestRequest_valid_1;
  wire                _zz_targets_0_bestRequest_priority_6;
  reg        [1:0]    targets_0_bestRequest_priority;
  reg        [4:0]    targets_0_bestRequest_id;
  reg                 targets_0_bestRequest_valid;
  wire                targets_0_iep;
  wire       [4:0]    targets_0_claim;
  wire                targets_1_ie_0;
  wire                targets_1_ie_1;
  wire                targets_1_ie_2;
  wire                targets_1_ie_3;
  wire                targets_1_ie_4;
  wire                targets_1_ie_5;
  wire                targets_1_ie_6;
  wire                targets_1_ie_7;
  wire                targets_1_ie_8;
  wire                targets_1_ie_9;
  wire                targets_1_ie_10;
  wire                targets_1_ie_11;
  wire                targets_1_ie_12;
  wire                targets_1_ie_13;
  wire                targets_1_ie_14;
  wire                targets_1_ie_15;
  wire                targets_1_ie_16;
  wire                targets_1_ie_17;
  wire                targets_1_ie_18;
  wire                targets_1_ie_19;
  wire                targets_1_ie_20;
  wire                targets_1_ie_21;
  wire                targets_1_ie_22;
  wire                targets_1_ie_23;
  wire                targets_1_ie_24;
  wire                targets_1_ie_25;
  wire                targets_1_ie_26;
  wire                targets_1_ie_27;
  wire                targets_1_ie_28;
  wire                targets_1_ie_29;
  wire                targets_1_ie_30;
  wire       [1:0]    targets_1_threshold;
  wire       [1:0]    targets_1_requests_0_priority;
  wire       [4:0]    targets_1_requests_0_id;
  wire                targets_1_requests_0_valid;
  wire       [1:0]    targets_1_requests_1_priority;
  wire       [4:0]    targets_1_requests_1_id;
  wire                targets_1_requests_1_valid;
  wire       [1:0]    targets_1_requests_2_priority;
  wire       [4:0]    targets_1_requests_2_id;
  wire                targets_1_requests_2_valid;
  wire       [1:0]    targets_1_requests_3_priority;
  wire       [4:0]    targets_1_requests_3_id;
  wire                targets_1_requests_3_valid;
  wire       [1:0]    targets_1_requests_4_priority;
  wire       [4:0]    targets_1_requests_4_id;
  wire                targets_1_requests_4_valid;
  wire       [1:0]    targets_1_requests_5_priority;
  wire       [4:0]    targets_1_requests_5_id;
  wire                targets_1_requests_5_valid;
  wire       [1:0]    targets_1_requests_6_priority;
  wire       [4:0]    targets_1_requests_6_id;
  wire                targets_1_requests_6_valid;
  wire       [1:0]    targets_1_requests_7_priority;
  wire       [4:0]    targets_1_requests_7_id;
  wire                targets_1_requests_7_valid;
  wire       [1:0]    targets_1_requests_8_priority;
  wire       [4:0]    targets_1_requests_8_id;
  wire                targets_1_requests_8_valid;
  wire       [1:0]    targets_1_requests_9_priority;
  wire       [4:0]    targets_1_requests_9_id;
  wire                targets_1_requests_9_valid;
  wire       [1:0]    targets_1_requests_10_priority;
  wire       [4:0]    targets_1_requests_10_id;
  wire                targets_1_requests_10_valid;
  wire       [1:0]    targets_1_requests_11_priority;
  wire       [4:0]    targets_1_requests_11_id;
  wire                targets_1_requests_11_valid;
  wire       [1:0]    targets_1_requests_12_priority;
  wire       [4:0]    targets_1_requests_12_id;
  wire                targets_1_requests_12_valid;
  wire       [1:0]    targets_1_requests_13_priority;
  wire       [4:0]    targets_1_requests_13_id;
  wire                targets_1_requests_13_valid;
  wire       [1:0]    targets_1_requests_14_priority;
  wire       [4:0]    targets_1_requests_14_id;
  wire                targets_1_requests_14_valid;
  wire       [1:0]    targets_1_requests_15_priority;
  wire       [4:0]    targets_1_requests_15_id;
  wire                targets_1_requests_15_valid;
  wire       [1:0]    targets_1_requests_16_priority;
  wire       [4:0]    targets_1_requests_16_id;
  wire                targets_1_requests_16_valid;
  wire       [1:0]    targets_1_requests_17_priority;
  wire       [4:0]    targets_1_requests_17_id;
  wire                targets_1_requests_17_valid;
  wire       [1:0]    targets_1_requests_18_priority;
  wire       [4:0]    targets_1_requests_18_id;
  wire                targets_1_requests_18_valid;
  wire       [1:0]    targets_1_requests_19_priority;
  wire       [4:0]    targets_1_requests_19_id;
  wire                targets_1_requests_19_valid;
  wire       [1:0]    targets_1_requests_20_priority;
  wire       [4:0]    targets_1_requests_20_id;
  wire                targets_1_requests_20_valid;
  wire       [1:0]    targets_1_requests_21_priority;
  wire       [4:0]    targets_1_requests_21_id;
  wire                targets_1_requests_21_valid;
  wire       [1:0]    targets_1_requests_22_priority;
  wire       [4:0]    targets_1_requests_22_id;
  wire                targets_1_requests_22_valid;
  wire       [1:0]    targets_1_requests_23_priority;
  wire       [4:0]    targets_1_requests_23_id;
  wire                targets_1_requests_23_valid;
  wire       [1:0]    targets_1_requests_24_priority;
  wire       [4:0]    targets_1_requests_24_id;
  wire                targets_1_requests_24_valid;
  wire       [1:0]    targets_1_requests_25_priority;
  wire       [4:0]    targets_1_requests_25_id;
  wire                targets_1_requests_25_valid;
  wire       [1:0]    targets_1_requests_26_priority;
  wire       [4:0]    targets_1_requests_26_id;
  wire                targets_1_requests_26_valid;
  wire       [1:0]    targets_1_requests_27_priority;
  wire       [4:0]    targets_1_requests_27_id;
  wire                targets_1_requests_27_valid;
  wire       [1:0]    targets_1_requests_28_priority;
  wire       [4:0]    targets_1_requests_28_id;
  wire                targets_1_requests_28_valid;
  wire       [1:0]    targets_1_requests_29_priority;
  wire       [4:0]    targets_1_requests_29_id;
  wire                targets_1_requests_29_valid;
  wire       [1:0]    targets_1_requests_30_priority;
  wire       [4:0]    targets_1_requests_30_id;
  wire                targets_1_requests_30_valid;
  wire       [1:0]    targets_1_requests_31_priority;
  wire       [4:0]    targets_1_requests_31_id;
  wire                targets_1_requests_31_valid;
  wire                _zz_targets_1_bestRequest_id;
  wire       [1:0]    _zz_targets_1_bestRequest_id_1;
  wire                _zz_targets_1_bestRequest_id_2;
  wire                _zz_targets_1_bestRequest_id_3;
  wire       [1:0]    _zz_targets_1_bestRequest_id_4;
  wire                _zz_targets_1_bestRequest_id_5;
  wire                _zz_targets_1_bestRequest_id_6;
  wire       [1:0]    _zz_targets_1_bestRequest_id_7;
  wire                _zz_targets_1_bestRequest_id_8;
  wire                _zz_targets_1_bestRequest_id_9;
  wire       [1:0]    _zz_targets_1_bestRequest_id_10;
  wire                _zz_targets_1_bestRequest_id_11;
  wire                _zz_targets_1_bestRequest_id_12;
  wire       [1:0]    _zz_targets_1_bestRequest_id_13;
  wire                _zz_targets_1_bestRequest_id_14;
  wire                _zz_targets_1_bestRequest_id_15;
  wire       [1:0]    _zz_targets_1_bestRequest_id_16;
  wire                _zz_targets_1_bestRequest_id_17;
  wire                _zz_targets_1_bestRequest_id_18;
  wire       [1:0]    _zz_targets_1_bestRequest_id_19;
  wire                _zz_targets_1_bestRequest_id_20;
  wire                _zz_targets_1_bestRequest_id_21;
  wire       [1:0]    _zz_targets_1_bestRequest_id_22;
  wire                _zz_targets_1_bestRequest_id_23;
  wire                _zz_targets_1_bestRequest_id_24;
  wire       [1:0]    _zz_targets_1_bestRequest_id_25;
  wire                _zz_targets_1_bestRequest_id_26;
  wire                _zz_targets_1_bestRequest_id_27;
  wire       [1:0]    _zz_targets_1_bestRequest_id_28;
  wire                _zz_targets_1_bestRequest_id_29;
  wire                _zz_targets_1_bestRequest_id_30;
  wire       [1:0]    _zz_targets_1_bestRequest_id_31;
  wire                _zz_targets_1_bestRequest_id_32;
  wire                _zz_targets_1_bestRequest_id_33;
  wire       [1:0]    _zz_targets_1_bestRequest_id_34;
  wire                _zz_targets_1_bestRequest_id_35;
  wire                _zz_targets_1_bestRequest_id_36;
  wire       [1:0]    _zz_targets_1_bestRequest_id_37;
  wire                _zz_targets_1_bestRequest_id_38;
  wire                _zz_targets_1_bestRequest_id_39;
  wire       [1:0]    _zz_targets_1_bestRequest_id_40;
  wire                _zz_targets_1_bestRequest_id_41;
  wire                _zz_targets_1_bestRequest_id_42;
  wire       [1:0]    _zz_targets_1_bestRequest_id_43;
  wire                _zz_targets_1_bestRequest_id_44;
  wire                _zz_targets_1_bestRequest_id_45;
  wire       [1:0]    _zz_targets_1_bestRequest_id_46;
  wire                _zz_targets_1_bestRequest_id_47;
  wire                _zz_targets_1_bestRequest_id_48;
  wire       [1:0]    _zz_targets_1_bestRequest_id_49;
  wire                _zz_targets_1_bestRequest_id_50;
  wire                _zz_targets_1_bestRequest_id_51;
  wire       [1:0]    _zz_targets_1_bestRequest_id_52;
  wire                _zz_targets_1_bestRequest_id_53;
  wire                _zz_targets_1_bestRequest_id_54;
  wire       [1:0]    _zz_targets_1_bestRequest_id_55;
  wire                _zz_targets_1_bestRequest_id_56;
  wire                _zz_targets_1_bestRequest_id_57;
  wire       [1:0]    _zz_targets_1_bestRequest_id_58;
  wire                _zz_targets_1_bestRequest_id_59;
  wire                _zz_targets_1_bestRequest_id_60;
  wire       [1:0]    _zz_targets_1_bestRequest_id_61;
  wire                _zz_targets_1_bestRequest_id_62;
  wire                _zz_targets_1_bestRequest_id_63;
  wire       [1:0]    _zz_targets_1_bestRequest_id_64;
  wire                _zz_targets_1_bestRequest_id_65;
  wire                _zz_targets_1_bestRequest_id_66;
  wire       [1:0]    _zz_targets_1_bestRequest_id_67;
  wire                _zz_targets_1_bestRequest_id_68;
  wire                _zz_targets_1_bestRequest_id_69;
  wire       [1:0]    _zz_targets_1_bestRequest_id_70;
  wire                _zz_targets_1_bestRequest_id_71;
  wire                _zz_targets_1_bestRequest_id_72;
  wire       [1:0]    _zz_targets_1_bestRequest_priority;
  wire                _zz_targets_1_bestRequest_id_73;
  wire                _zz_targets_1_bestRequest_id_74;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_1;
  wire                _zz_targets_1_bestRequest_id_75;
  wire                _zz_targets_1_bestRequest_id_76;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_2;
  wire                _zz_targets_1_bestRequest_id_77;
  wire                _zz_targets_1_bestRequest_id_78;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_3;
  wire                _zz_targets_1_bestRequest_id_79;
  wire                _zz_targets_1_bestRequest_id_80;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_4;
  wire                _zz_targets_1_bestRequest_valid;
  wire                _zz_targets_1_bestRequest_id_81;
  wire       [1:0]    _zz_targets_1_bestRequest_priority_5;
  wire                _zz_targets_1_bestRequest_valid_1;
  wire                _zz_targets_1_bestRequest_priority_6;
  reg        [1:0]    targets_1_bestRequest_priority;
  reg        [4:0]    targets_1_bestRequest_id;
  reg                 targets_1_bestRequest_valid;
  wire                targets_1_iep;
  wire       [4:0]    targets_1_claim;
  wire                factory_readErrorFlag;
  wire                factory_writeErrorFlag;
  wire                factory_rspAsync_valid;
  reg                 factory_rspAsync_ready;
  wire       [2:0]    factory_rspAsync_payload_opcode;
  wire       [2:0]    factory_rspAsync_payload_param;
  wire       [2:0]    factory_rspAsync_payload_source;
  wire       [1:0]    factory_rspAsync_payload_size;
  wire                factory_rspAsync_payload_denied;
  reg        [31:0]   factory_rspAsync_payload_data;
  wire                factory_rspAsync_payload_corrupt;
  wire                factory_askWrite;
  wire                factory_askRead;
  wire                factory_doWrite;
  wire                factory_doRead;
  wire       [21:0]   factory_address;
  reg                 factory_halt;
  reg        [1:0]    gateways_0_priority_driver;
  reg        [1:0]    gateways_1_priority_driver;
  reg        [1:0]    gateways_2_priority_driver;
  reg        [1:0]    gateways_3_priority_driver;
  reg        [1:0]    gateways_4_priority_driver;
  reg        [1:0]    gateways_5_priority_driver;
  reg        [1:0]    gateways_6_priority_driver;
  reg        [1:0]    gateways_7_priority_driver;
  reg        [1:0]    gateways_8_priority_driver;
  reg        [1:0]    gateways_9_priority_driver;
  reg        [1:0]    gateways_10_priority_driver;
  reg        [1:0]    gateways_11_priority_driver;
  reg        [1:0]    gateways_12_priority_driver;
  reg        [1:0]    gateways_13_priority_driver;
  reg        [1:0]    gateways_14_priority_driver;
  reg        [1:0]    gateways_15_priority_driver;
  reg        [1:0]    gateways_16_priority_driver;
  reg        [1:0]    gateways_17_priority_driver;
  reg        [1:0]    gateways_18_priority_driver;
  reg        [1:0]    gateways_19_priority_driver;
  reg        [1:0]    gateways_20_priority_driver;
  reg        [1:0]    gateways_21_priority_driver;
  reg        [1:0]    gateways_22_priority_driver;
  reg        [1:0]    gateways_23_priority_driver;
  reg        [1:0]    gateways_24_priority_driver;
  reg        [1:0]    gateways_25_priority_driver;
  reg        [1:0]    gateways_26_priority_driver;
  reg        [1:0]    gateways_27_priority_driver;
  reg        [1:0]    gateways_28_priority_driver;
  reg        [1:0]    gateways_29_priority_driver;
  reg        [1:0]    gateways_30_priority_driver;
  reg                 mapping_claim_valid;
  reg        [4:0]    mapping_claim_payload;
  reg                 mapping_completion_valid;
  reg        [4:0]    mapping_completion_payload;
  reg                 mapping_coherencyStall_willIncrement;
  wire                mapping_coherencyStall_willClear;
  reg        [0:0]    mapping_coherencyStall_valueNext;
  reg        [0:0]    mapping_coherencyStall_value;
  wire                mapping_coherencyStall_willOverflowIfInc;
  wire                mapping_coherencyStall_willOverflow;
  wire                when_PlicMapper_l122;
  reg        [1:0]    targets_0_threshold_driver;
  reg                 mapping_targetMapping_0_targetCompletion_valid;
  wire       [4:0]    mapping_targetMapping_0_targetCompletion_payload;
  reg                 targets_0_ie_0_driver;
  reg                 targets_0_ie_1_driver;
  reg                 targets_0_ie_2_driver;
  reg                 targets_0_ie_3_driver;
  reg                 targets_0_ie_4_driver;
  reg                 targets_0_ie_5_driver;
  reg                 targets_0_ie_6_driver;
  reg                 targets_0_ie_7_driver;
  reg                 targets_0_ie_8_driver;
  reg                 targets_0_ie_9_driver;
  reg                 targets_0_ie_10_driver;
  reg                 targets_0_ie_11_driver;
  reg                 targets_0_ie_12_driver;
  reg                 targets_0_ie_13_driver;
  reg                 targets_0_ie_14_driver;
  reg                 targets_0_ie_15_driver;
  reg                 targets_0_ie_16_driver;
  reg                 targets_0_ie_17_driver;
  reg                 targets_0_ie_18_driver;
  reg                 targets_0_ie_19_driver;
  reg                 targets_0_ie_20_driver;
  reg                 targets_0_ie_21_driver;
  reg                 targets_0_ie_22_driver;
  reg                 targets_0_ie_23_driver;
  reg                 targets_0_ie_24_driver;
  reg                 targets_0_ie_25_driver;
  reg                 targets_0_ie_26_driver;
  reg                 targets_0_ie_27_driver;
  reg                 targets_0_ie_28_driver;
  reg                 targets_0_ie_29_driver;
  reg                 targets_0_ie_30_driver;
  reg        [1:0]    targets_1_threshold_driver;
  reg                 mapping_targetMapping_1_targetCompletion_valid;
  wire       [4:0]    mapping_targetMapping_1_targetCompletion_payload;
  reg                 targets_1_ie_0_driver;
  reg                 targets_1_ie_1_driver;
  reg                 targets_1_ie_2_driver;
  reg                 targets_1_ie_3_driver;
  reg                 targets_1_ie_4_driver;
  reg                 targets_1_ie_5_driver;
  reg                 targets_1_ie_6_driver;
  reg                 targets_1_ie_7_driver;
  reg                 targets_1_ie_8_driver;
  reg                 targets_1_ie_9_driver;
  reg                 targets_1_ie_10_driver;
  reg                 targets_1_ie_11_driver;
  reg                 targets_1_ie_12_driver;
  reg                 targets_1_ie_13_driver;
  reg                 targets_1_ie_14_driver;
  reg                 targets_1_ie_15_driver;
  reg                 targets_1_ie_16_driver;
  reg                 targets_1_ie_17_driver;
  reg                 targets_1_ie_18_driver;
  reg                 targets_1_ie_19_driver;
  reg                 targets_1_ie_20_driver;
  reg                 targets_1_ie_21_driver;
  reg                 targets_1_ie_22_driver;
  reg                 targets_1_ie_23_driver;
  reg                 targets_1_ie_24_driver;
  reg                 targets_1_ie_25_driver;
  reg                 targets_1_ie_26_driver;
  reg                 targets_1_ie_27_driver;
  reg                 targets_1_ie_28_driver;
  reg                 targets_1_ie_29_driver;
  reg                 targets_1_ie_30_driver;
  wire       [2:0]    _zz_factory_rspAsync_payload_opcode;
  wire                factory_rspAsync_stage_valid;
  wire                factory_rspAsync_stage_ready;
  wire       [2:0]    factory_rspAsync_stage_payload_opcode;
  wire       [2:0]    factory_rspAsync_stage_payload_param;
  wire       [2:0]    factory_rspAsync_stage_payload_source;
  wire       [1:0]    factory_rspAsync_stage_payload_size;
  wire                factory_rspAsync_stage_payload_denied;
  wire       [31:0]   factory_rspAsync_stage_payload_data;
  wire                factory_rspAsync_stage_payload_corrupt;
  reg                 factory_rspAsync_rValid;
  reg        [2:0]    factory_rspAsync_rData_opcode;
  reg        [2:0]    factory_rspAsync_rData_param;
  reg        [2:0]    factory_rspAsync_rData_source;
  reg        [1:0]    factory_rspAsync_rData_size;
  reg                 factory_rspAsync_rData_denied;
  reg        [31:0]   factory_rspAsync_rData_data;
  reg                 factory_rspAsync_rData_corrupt;
  wire                when_Stream_l399;
  wire                when_SlaveFactory_l134;
  `ifndef SYNTHESIS
  reg [127:0] io_bus_a_payload_opcode_string;
  reg [119:0] io_bus_d_payload_opcode_string;
  reg [119:0] factory_rspAsync_payload_opcode_string;
  reg [119:0] _zz_factory_rspAsync_payload_opcode_string;
  reg [119:0] factory_rspAsync_stage_payload_opcode_string;
  reg [119:0] factory_rspAsync_rData_opcode_string;
  `endif


  assign _zz_factory_address = (io_bus_a_payload_address >>> 2'd2);
  assign _zz_targets_0_bestRequest_id_82 = (_zz_targets_0_bestRequest_id ? targets_0_requests_0_id : targets_0_requests_1_id);
  assign _zz_targets_0_bestRequest_id_83 = (_zz_targets_0_bestRequest_id_3 ? targets_0_requests_2_id : targets_0_requests_3_id);
  assign _zz_targets_0_bestRequest_id_84 = (_zz_targets_0_bestRequest_id_6 ? targets_0_requests_4_id : targets_0_requests_5_id);
  assign _zz_targets_0_bestRequest_id_85 = (_zz_targets_0_bestRequest_id_9 ? targets_0_requests_6_id : targets_0_requests_7_id);
  assign _zz_targets_0_bestRequest_id_86 = (_zz_targets_0_bestRequest_id_12 ? targets_0_requests_8_id : targets_0_requests_9_id);
  assign _zz_targets_0_bestRequest_id_87 = (_zz_targets_0_bestRequest_id_15 ? targets_0_requests_10_id : targets_0_requests_11_id);
  assign _zz_targets_0_bestRequest_id_88 = (_zz_targets_0_bestRequest_id_18 ? targets_0_requests_12_id : targets_0_requests_13_id);
  assign _zz_targets_0_bestRequest_id_89 = (_zz_targets_0_bestRequest_id_21 ? targets_0_requests_14_id : targets_0_requests_15_id);
  assign _zz_targets_0_bestRequest_id_90 = (_zz_targets_0_bestRequest_id_24 ? targets_0_requests_16_id : targets_0_requests_17_id);
  assign _zz_targets_0_bestRequest_id_91 = (_zz_targets_0_bestRequest_id_27 ? targets_0_requests_18_id : targets_0_requests_19_id);
  assign _zz_targets_0_bestRequest_id_92 = (_zz_targets_0_bestRequest_id_30 ? targets_0_requests_20_id : targets_0_requests_21_id);
  assign _zz_targets_0_bestRequest_id_93 = (_zz_targets_0_bestRequest_id_33 ? targets_0_requests_22_id : targets_0_requests_23_id);
  assign _zz_targets_0_bestRequest_id_94 = (_zz_targets_0_bestRequest_id_36 ? targets_0_requests_24_id : targets_0_requests_25_id);
  assign _zz_targets_0_bestRequest_id_95 = (_zz_targets_0_bestRequest_id_39 ? targets_0_requests_26_id : targets_0_requests_27_id);
  assign _zz_targets_0_bestRequest_id_96 = (_zz_targets_0_bestRequest_id_42 ? targets_0_requests_28_id : targets_0_requests_29_id);
  assign _zz_targets_0_bestRequest_id_97 = (_zz_targets_0_bestRequest_id_45 ? targets_0_requests_30_id : targets_0_requests_31_id);
  assign _zz_targets_1_bestRequest_id_82 = (_zz_targets_1_bestRequest_id ? targets_1_requests_0_id : targets_1_requests_1_id);
  assign _zz_targets_1_bestRequest_id_83 = (_zz_targets_1_bestRequest_id_3 ? targets_1_requests_2_id : targets_1_requests_3_id);
  assign _zz_targets_1_bestRequest_id_84 = (_zz_targets_1_bestRequest_id_6 ? targets_1_requests_4_id : targets_1_requests_5_id);
  assign _zz_targets_1_bestRequest_id_85 = (_zz_targets_1_bestRequest_id_9 ? targets_1_requests_6_id : targets_1_requests_7_id);
  assign _zz_targets_1_bestRequest_id_86 = (_zz_targets_1_bestRequest_id_12 ? targets_1_requests_8_id : targets_1_requests_9_id);
  assign _zz_targets_1_bestRequest_id_87 = (_zz_targets_1_bestRequest_id_15 ? targets_1_requests_10_id : targets_1_requests_11_id);
  assign _zz_targets_1_bestRequest_id_88 = (_zz_targets_1_bestRequest_id_18 ? targets_1_requests_12_id : targets_1_requests_13_id);
  assign _zz_targets_1_bestRequest_id_89 = (_zz_targets_1_bestRequest_id_21 ? targets_1_requests_14_id : targets_1_requests_15_id);
  assign _zz_targets_1_bestRequest_id_90 = (_zz_targets_1_bestRequest_id_24 ? targets_1_requests_16_id : targets_1_requests_17_id);
  assign _zz_targets_1_bestRequest_id_91 = (_zz_targets_1_bestRequest_id_27 ? targets_1_requests_18_id : targets_1_requests_19_id);
  assign _zz_targets_1_bestRequest_id_92 = (_zz_targets_1_bestRequest_id_30 ? targets_1_requests_20_id : targets_1_requests_21_id);
  assign _zz_targets_1_bestRequest_id_93 = (_zz_targets_1_bestRequest_id_33 ? targets_1_requests_22_id : targets_1_requests_23_id);
  assign _zz_targets_1_bestRequest_id_94 = (_zz_targets_1_bestRequest_id_36 ? targets_1_requests_24_id : targets_1_requests_25_id);
  assign _zz_targets_1_bestRequest_id_95 = (_zz_targets_1_bestRequest_id_39 ? targets_1_requests_26_id : targets_1_requests_27_id);
  assign _zz_targets_1_bestRequest_id_96 = (_zz_targets_1_bestRequest_id_42 ? targets_1_requests_28_id : targets_1_requests_29_id);
  assign _zz_targets_1_bestRequest_id_97 = (_zz_targets_1_bestRequest_id_45 ? targets_1_requests_30_id : targets_1_requests_31_id);
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_bus_a_payload_opcode)
      A_PUT_FULL_DATA : io_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_bus_d_payload_opcode)
      D_ACCESS_ACK : io_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(factory_rspAsync_payload_opcode)
      D_ACCESS_ACK : factory_rspAsync_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : factory_rspAsync_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : factory_rspAsync_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : factory_rspAsync_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : factory_rspAsync_payload_opcode_string = "RELEASE_ACK    ";
      default : factory_rspAsync_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_factory_rspAsync_payload_opcode)
      D_ACCESS_ACK : _zz_factory_rspAsync_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_factory_rspAsync_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_factory_rspAsync_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_factory_rspAsync_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_factory_rspAsync_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_factory_rspAsync_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(factory_rspAsync_stage_payload_opcode)
      D_ACCESS_ACK : factory_rspAsync_stage_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : factory_rspAsync_stage_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : factory_rspAsync_stage_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : factory_rspAsync_stage_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : factory_rspAsync_stage_payload_opcode_string = "RELEASE_ACK    ";
      default : factory_rspAsync_stage_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(factory_rspAsync_rData_opcode)
      D_ACCESS_ACK : factory_rspAsync_rData_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : factory_rspAsync_rData_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : factory_rspAsync_rData_opcode_string = "GRANT          ";
      D_GRANT_DATA : factory_rspAsync_rData_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : factory_rspAsync_rData_opcode_string = "RELEASE_ACK    ";
      default : factory_rspAsync_rData_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign _zz_gateways_0_ip = io_sources[0];
  assign _zz_gateways_1_ip = io_sources[1];
  assign _zz_gateways_2_ip = io_sources[2];
  assign _zz_gateways_3_ip = io_sources[3];
  assign _zz_gateways_4_ip = io_sources[4];
  assign _zz_gateways_5_ip = io_sources[5];
  assign _zz_gateways_6_ip = io_sources[6];
  assign _zz_gateways_7_ip = io_sources[7];
  assign _zz_gateways_8_ip = io_sources[8];
  assign _zz_gateways_9_ip = io_sources[9];
  assign _zz_gateways_10_ip = io_sources[10];
  assign _zz_gateways_11_ip = io_sources[11];
  assign _zz_gateways_12_ip = io_sources[12];
  assign _zz_gateways_13_ip = io_sources[13];
  assign _zz_gateways_14_ip = io_sources[14];
  assign _zz_gateways_15_ip = io_sources[15];
  assign _zz_gateways_16_ip = io_sources[16];
  assign _zz_gateways_17_ip = io_sources[17];
  assign _zz_gateways_18_ip = io_sources[18];
  assign _zz_gateways_19_ip = io_sources[19];
  assign _zz_gateways_20_ip = io_sources[20];
  assign _zz_gateways_21_ip = io_sources[21];
  assign _zz_gateways_22_ip = io_sources[22];
  assign _zz_gateways_23_ip = io_sources[23];
  assign _zz_gateways_24_ip = io_sources[24];
  assign _zz_gateways_25_ip = io_sources[25];
  assign _zz_gateways_26_ip = io_sources[26];
  assign _zz_gateways_27_ip = io_sources[27];
  assign _zz_gateways_28_ip = io_sources[28];
  assign _zz_gateways_29_ip = io_sources[29];
  assign _zz_gateways_30_ip = io_sources[30];
  assign when_PlicGateway_l21 = (! gateways_0_waitCompletion);
  assign when_PlicGateway_l21_1 = (! gateways_1_waitCompletion);
  assign when_PlicGateway_l21_2 = (! gateways_2_waitCompletion);
  assign when_PlicGateway_l21_3 = (! gateways_3_waitCompletion);
  assign when_PlicGateway_l21_4 = (! gateways_4_waitCompletion);
  assign when_PlicGateway_l21_5 = (! gateways_5_waitCompletion);
  assign when_PlicGateway_l21_6 = (! gateways_6_waitCompletion);
  assign when_PlicGateway_l21_7 = (! gateways_7_waitCompletion);
  assign when_PlicGateway_l21_8 = (! gateways_8_waitCompletion);
  assign when_PlicGateway_l21_9 = (! gateways_9_waitCompletion);
  assign when_PlicGateway_l21_10 = (! gateways_10_waitCompletion);
  assign when_PlicGateway_l21_11 = (! gateways_11_waitCompletion);
  assign when_PlicGateway_l21_12 = (! gateways_12_waitCompletion);
  assign when_PlicGateway_l21_13 = (! gateways_13_waitCompletion);
  assign when_PlicGateway_l21_14 = (! gateways_14_waitCompletion);
  assign when_PlicGateway_l21_15 = (! gateways_15_waitCompletion);
  assign when_PlicGateway_l21_16 = (! gateways_16_waitCompletion);
  assign when_PlicGateway_l21_17 = (! gateways_17_waitCompletion);
  assign when_PlicGateway_l21_18 = (! gateways_18_waitCompletion);
  assign when_PlicGateway_l21_19 = (! gateways_19_waitCompletion);
  assign when_PlicGateway_l21_20 = (! gateways_20_waitCompletion);
  assign when_PlicGateway_l21_21 = (! gateways_21_waitCompletion);
  assign when_PlicGateway_l21_22 = (! gateways_22_waitCompletion);
  assign when_PlicGateway_l21_23 = (! gateways_23_waitCompletion);
  assign when_PlicGateway_l21_24 = (! gateways_24_waitCompletion);
  assign when_PlicGateway_l21_25 = (! gateways_25_waitCompletion);
  assign when_PlicGateway_l21_26 = (! gateways_26_waitCompletion);
  assign when_PlicGateway_l21_27 = (! gateways_27_waitCompletion);
  assign when_PlicGateway_l21_28 = (! gateways_28_waitCompletion);
  assign when_PlicGateway_l21_29 = (! gateways_29_waitCompletion);
  assign when_PlicGateway_l21_30 = (! gateways_30_waitCompletion);
  assign targets_0_requests_0_priority = 2'b00;
  assign targets_0_requests_0_id = 5'h0;
  assign targets_0_requests_0_valid = 1'b1;
  assign targets_0_requests_1_priority = gateways_0_priority;
  assign targets_0_requests_1_id = 5'h01;
  assign targets_0_requests_1_valid = (gateways_0_ip && targets_0_ie_0);
  assign targets_0_requests_2_priority = gateways_1_priority;
  assign targets_0_requests_2_id = 5'h02;
  assign targets_0_requests_2_valid = (gateways_1_ip && targets_0_ie_1);
  assign targets_0_requests_3_priority = gateways_2_priority;
  assign targets_0_requests_3_id = 5'h03;
  assign targets_0_requests_3_valid = (gateways_2_ip && targets_0_ie_2);
  assign targets_0_requests_4_priority = gateways_3_priority;
  assign targets_0_requests_4_id = 5'h04;
  assign targets_0_requests_4_valid = (gateways_3_ip && targets_0_ie_3);
  assign targets_0_requests_5_priority = gateways_4_priority;
  assign targets_0_requests_5_id = 5'h05;
  assign targets_0_requests_5_valid = (gateways_4_ip && targets_0_ie_4);
  assign targets_0_requests_6_priority = gateways_5_priority;
  assign targets_0_requests_6_id = 5'h06;
  assign targets_0_requests_6_valid = (gateways_5_ip && targets_0_ie_5);
  assign targets_0_requests_7_priority = gateways_6_priority;
  assign targets_0_requests_7_id = 5'h07;
  assign targets_0_requests_7_valid = (gateways_6_ip && targets_0_ie_6);
  assign targets_0_requests_8_priority = gateways_7_priority;
  assign targets_0_requests_8_id = 5'h08;
  assign targets_0_requests_8_valid = (gateways_7_ip && targets_0_ie_7);
  assign targets_0_requests_9_priority = gateways_8_priority;
  assign targets_0_requests_9_id = 5'h09;
  assign targets_0_requests_9_valid = (gateways_8_ip && targets_0_ie_8);
  assign targets_0_requests_10_priority = gateways_9_priority;
  assign targets_0_requests_10_id = 5'h0a;
  assign targets_0_requests_10_valid = (gateways_9_ip && targets_0_ie_9);
  assign targets_0_requests_11_priority = gateways_10_priority;
  assign targets_0_requests_11_id = 5'h0b;
  assign targets_0_requests_11_valid = (gateways_10_ip && targets_0_ie_10);
  assign targets_0_requests_12_priority = gateways_11_priority;
  assign targets_0_requests_12_id = 5'h0c;
  assign targets_0_requests_12_valid = (gateways_11_ip && targets_0_ie_11);
  assign targets_0_requests_13_priority = gateways_12_priority;
  assign targets_0_requests_13_id = 5'h0d;
  assign targets_0_requests_13_valid = (gateways_12_ip && targets_0_ie_12);
  assign targets_0_requests_14_priority = gateways_13_priority;
  assign targets_0_requests_14_id = 5'h0e;
  assign targets_0_requests_14_valid = (gateways_13_ip && targets_0_ie_13);
  assign targets_0_requests_15_priority = gateways_14_priority;
  assign targets_0_requests_15_id = 5'h0f;
  assign targets_0_requests_15_valid = (gateways_14_ip && targets_0_ie_14);
  assign targets_0_requests_16_priority = gateways_15_priority;
  assign targets_0_requests_16_id = 5'h10;
  assign targets_0_requests_16_valid = (gateways_15_ip && targets_0_ie_15);
  assign targets_0_requests_17_priority = gateways_16_priority;
  assign targets_0_requests_17_id = 5'h11;
  assign targets_0_requests_17_valid = (gateways_16_ip && targets_0_ie_16);
  assign targets_0_requests_18_priority = gateways_17_priority;
  assign targets_0_requests_18_id = 5'h12;
  assign targets_0_requests_18_valid = (gateways_17_ip && targets_0_ie_17);
  assign targets_0_requests_19_priority = gateways_18_priority;
  assign targets_0_requests_19_id = 5'h13;
  assign targets_0_requests_19_valid = (gateways_18_ip && targets_0_ie_18);
  assign targets_0_requests_20_priority = gateways_19_priority;
  assign targets_0_requests_20_id = 5'h14;
  assign targets_0_requests_20_valid = (gateways_19_ip && targets_0_ie_19);
  assign targets_0_requests_21_priority = gateways_20_priority;
  assign targets_0_requests_21_id = 5'h15;
  assign targets_0_requests_21_valid = (gateways_20_ip && targets_0_ie_20);
  assign targets_0_requests_22_priority = gateways_21_priority;
  assign targets_0_requests_22_id = 5'h16;
  assign targets_0_requests_22_valid = (gateways_21_ip && targets_0_ie_21);
  assign targets_0_requests_23_priority = gateways_22_priority;
  assign targets_0_requests_23_id = 5'h17;
  assign targets_0_requests_23_valid = (gateways_22_ip && targets_0_ie_22);
  assign targets_0_requests_24_priority = gateways_23_priority;
  assign targets_0_requests_24_id = 5'h18;
  assign targets_0_requests_24_valid = (gateways_23_ip && targets_0_ie_23);
  assign targets_0_requests_25_priority = gateways_24_priority;
  assign targets_0_requests_25_id = 5'h19;
  assign targets_0_requests_25_valid = (gateways_24_ip && targets_0_ie_24);
  assign targets_0_requests_26_priority = gateways_25_priority;
  assign targets_0_requests_26_id = 5'h1a;
  assign targets_0_requests_26_valid = (gateways_25_ip && targets_0_ie_25);
  assign targets_0_requests_27_priority = gateways_26_priority;
  assign targets_0_requests_27_id = 5'h1b;
  assign targets_0_requests_27_valid = (gateways_26_ip && targets_0_ie_26);
  assign targets_0_requests_28_priority = gateways_27_priority;
  assign targets_0_requests_28_id = 5'h1c;
  assign targets_0_requests_28_valid = (gateways_27_ip && targets_0_ie_27);
  assign targets_0_requests_29_priority = gateways_28_priority;
  assign targets_0_requests_29_id = 5'h1d;
  assign targets_0_requests_29_valid = (gateways_28_ip && targets_0_ie_28);
  assign targets_0_requests_30_priority = gateways_29_priority;
  assign targets_0_requests_30_id = 5'h1e;
  assign targets_0_requests_30_valid = (gateways_29_ip && targets_0_ie_29);
  assign targets_0_requests_31_priority = gateways_30_priority;
  assign targets_0_requests_31_id = 5'h1f;
  assign targets_0_requests_31_valid = (gateways_30_ip && targets_0_ie_30);
  assign _zz_targets_0_bestRequest_id = ((! targets_0_requests_1_valid) || (targets_0_requests_0_valid && (targets_0_requests_1_priority <= targets_0_requests_0_priority)));
  assign _zz_targets_0_bestRequest_id_1 = (_zz_targets_0_bestRequest_id ? targets_0_requests_0_priority : targets_0_requests_1_priority);
  assign _zz_targets_0_bestRequest_id_2 = (_zz_targets_0_bestRequest_id ? targets_0_requests_0_valid : targets_0_requests_1_valid);
  assign _zz_targets_0_bestRequest_id_3 = ((! targets_0_requests_3_valid) || (targets_0_requests_2_valid && (targets_0_requests_3_priority <= targets_0_requests_2_priority)));
  assign _zz_targets_0_bestRequest_id_4 = (_zz_targets_0_bestRequest_id_3 ? targets_0_requests_2_priority : targets_0_requests_3_priority);
  assign _zz_targets_0_bestRequest_id_5 = (_zz_targets_0_bestRequest_id_3 ? targets_0_requests_2_valid : targets_0_requests_3_valid);
  assign _zz_targets_0_bestRequest_id_6 = ((! targets_0_requests_5_valid) || (targets_0_requests_4_valid && (targets_0_requests_5_priority <= targets_0_requests_4_priority)));
  assign _zz_targets_0_bestRequest_id_7 = (_zz_targets_0_bestRequest_id_6 ? targets_0_requests_4_priority : targets_0_requests_5_priority);
  assign _zz_targets_0_bestRequest_id_8 = (_zz_targets_0_bestRequest_id_6 ? targets_0_requests_4_valid : targets_0_requests_5_valid);
  assign _zz_targets_0_bestRequest_id_9 = ((! targets_0_requests_7_valid) || (targets_0_requests_6_valid && (targets_0_requests_7_priority <= targets_0_requests_6_priority)));
  assign _zz_targets_0_bestRequest_id_10 = (_zz_targets_0_bestRequest_id_9 ? targets_0_requests_6_priority : targets_0_requests_7_priority);
  assign _zz_targets_0_bestRequest_id_11 = (_zz_targets_0_bestRequest_id_9 ? targets_0_requests_6_valid : targets_0_requests_7_valid);
  assign _zz_targets_0_bestRequest_id_12 = ((! targets_0_requests_9_valid) || (targets_0_requests_8_valid && (targets_0_requests_9_priority <= targets_0_requests_8_priority)));
  assign _zz_targets_0_bestRequest_id_13 = (_zz_targets_0_bestRequest_id_12 ? targets_0_requests_8_priority : targets_0_requests_9_priority);
  assign _zz_targets_0_bestRequest_id_14 = (_zz_targets_0_bestRequest_id_12 ? targets_0_requests_8_valid : targets_0_requests_9_valid);
  assign _zz_targets_0_bestRequest_id_15 = ((! targets_0_requests_11_valid) || (targets_0_requests_10_valid && (targets_0_requests_11_priority <= targets_0_requests_10_priority)));
  assign _zz_targets_0_bestRequest_id_16 = (_zz_targets_0_bestRequest_id_15 ? targets_0_requests_10_priority : targets_0_requests_11_priority);
  assign _zz_targets_0_bestRequest_id_17 = (_zz_targets_0_bestRequest_id_15 ? targets_0_requests_10_valid : targets_0_requests_11_valid);
  assign _zz_targets_0_bestRequest_id_18 = ((! targets_0_requests_13_valid) || (targets_0_requests_12_valid && (targets_0_requests_13_priority <= targets_0_requests_12_priority)));
  assign _zz_targets_0_bestRequest_id_19 = (_zz_targets_0_bestRequest_id_18 ? targets_0_requests_12_priority : targets_0_requests_13_priority);
  assign _zz_targets_0_bestRequest_id_20 = (_zz_targets_0_bestRequest_id_18 ? targets_0_requests_12_valid : targets_0_requests_13_valid);
  assign _zz_targets_0_bestRequest_id_21 = ((! targets_0_requests_15_valid) || (targets_0_requests_14_valid && (targets_0_requests_15_priority <= targets_0_requests_14_priority)));
  assign _zz_targets_0_bestRequest_id_22 = (_zz_targets_0_bestRequest_id_21 ? targets_0_requests_14_priority : targets_0_requests_15_priority);
  assign _zz_targets_0_bestRequest_id_23 = (_zz_targets_0_bestRequest_id_21 ? targets_0_requests_14_valid : targets_0_requests_15_valid);
  assign _zz_targets_0_bestRequest_id_24 = ((! targets_0_requests_17_valid) || (targets_0_requests_16_valid && (targets_0_requests_17_priority <= targets_0_requests_16_priority)));
  assign _zz_targets_0_bestRequest_id_25 = (_zz_targets_0_bestRequest_id_24 ? targets_0_requests_16_priority : targets_0_requests_17_priority);
  assign _zz_targets_0_bestRequest_id_26 = (_zz_targets_0_bestRequest_id_24 ? targets_0_requests_16_valid : targets_0_requests_17_valid);
  assign _zz_targets_0_bestRequest_id_27 = ((! targets_0_requests_19_valid) || (targets_0_requests_18_valid && (targets_0_requests_19_priority <= targets_0_requests_18_priority)));
  assign _zz_targets_0_bestRequest_id_28 = (_zz_targets_0_bestRequest_id_27 ? targets_0_requests_18_priority : targets_0_requests_19_priority);
  assign _zz_targets_0_bestRequest_id_29 = (_zz_targets_0_bestRequest_id_27 ? targets_0_requests_18_valid : targets_0_requests_19_valid);
  assign _zz_targets_0_bestRequest_id_30 = ((! targets_0_requests_21_valid) || (targets_0_requests_20_valid && (targets_0_requests_21_priority <= targets_0_requests_20_priority)));
  assign _zz_targets_0_bestRequest_id_31 = (_zz_targets_0_bestRequest_id_30 ? targets_0_requests_20_priority : targets_0_requests_21_priority);
  assign _zz_targets_0_bestRequest_id_32 = (_zz_targets_0_bestRequest_id_30 ? targets_0_requests_20_valid : targets_0_requests_21_valid);
  assign _zz_targets_0_bestRequest_id_33 = ((! targets_0_requests_23_valid) || (targets_0_requests_22_valid && (targets_0_requests_23_priority <= targets_0_requests_22_priority)));
  assign _zz_targets_0_bestRequest_id_34 = (_zz_targets_0_bestRequest_id_33 ? targets_0_requests_22_priority : targets_0_requests_23_priority);
  assign _zz_targets_0_bestRequest_id_35 = (_zz_targets_0_bestRequest_id_33 ? targets_0_requests_22_valid : targets_0_requests_23_valid);
  assign _zz_targets_0_bestRequest_id_36 = ((! targets_0_requests_25_valid) || (targets_0_requests_24_valid && (targets_0_requests_25_priority <= targets_0_requests_24_priority)));
  assign _zz_targets_0_bestRequest_id_37 = (_zz_targets_0_bestRequest_id_36 ? targets_0_requests_24_priority : targets_0_requests_25_priority);
  assign _zz_targets_0_bestRequest_id_38 = (_zz_targets_0_bestRequest_id_36 ? targets_0_requests_24_valid : targets_0_requests_25_valid);
  assign _zz_targets_0_bestRequest_id_39 = ((! targets_0_requests_27_valid) || (targets_0_requests_26_valid && (targets_0_requests_27_priority <= targets_0_requests_26_priority)));
  assign _zz_targets_0_bestRequest_id_40 = (_zz_targets_0_bestRequest_id_39 ? targets_0_requests_26_priority : targets_0_requests_27_priority);
  assign _zz_targets_0_bestRequest_id_41 = (_zz_targets_0_bestRequest_id_39 ? targets_0_requests_26_valid : targets_0_requests_27_valid);
  assign _zz_targets_0_bestRequest_id_42 = ((! targets_0_requests_29_valid) || (targets_0_requests_28_valid && (targets_0_requests_29_priority <= targets_0_requests_28_priority)));
  assign _zz_targets_0_bestRequest_id_43 = (_zz_targets_0_bestRequest_id_42 ? targets_0_requests_28_priority : targets_0_requests_29_priority);
  assign _zz_targets_0_bestRequest_id_44 = (_zz_targets_0_bestRequest_id_42 ? targets_0_requests_28_valid : targets_0_requests_29_valid);
  assign _zz_targets_0_bestRequest_id_45 = ((! targets_0_requests_31_valid) || (targets_0_requests_30_valid && (targets_0_requests_31_priority <= targets_0_requests_30_priority)));
  assign _zz_targets_0_bestRequest_id_46 = (_zz_targets_0_bestRequest_id_45 ? targets_0_requests_30_priority : targets_0_requests_31_priority);
  assign _zz_targets_0_bestRequest_id_47 = (_zz_targets_0_bestRequest_id_45 ? targets_0_requests_30_valid : targets_0_requests_31_valid);
  assign _zz_targets_0_bestRequest_id_48 = ((! _zz_targets_0_bestRequest_id_5) || (_zz_targets_0_bestRequest_id_2 && (_zz_targets_0_bestRequest_id_4 <= _zz_targets_0_bestRequest_id_1)));
  assign _zz_targets_0_bestRequest_id_49 = (_zz_targets_0_bestRequest_id_48 ? _zz_targets_0_bestRequest_id_1 : _zz_targets_0_bestRequest_id_4);
  assign _zz_targets_0_bestRequest_id_50 = (_zz_targets_0_bestRequest_id_48 ? _zz_targets_0_bestRequest_id_2 : _zz_targets_0_bestRequest_id_5);
  assign _zz_targets_0_bestRequest_id_51 = ((! _zz_targets_0_bestRequest_id_11) || (_zz_targets_0_bestRequest_id_8 && (_zz_targets_0_bestRequest_id_10 <= _zz_targets_0_bestRequest_id_7)));
  assign _zz_targets_0_bestRequest_id_52 = (_zz_targets_0_bestRequest_id_51 ? _zz_targets_0_bestRequest_id_7 : _zz_targets_0_bestRequest_id_10);
  assign _zz_targets_0_bestRequest_id_53 = (_zz_targets_0_bestRequest_id_51 ? _zz_targets_0_bestRequest_id_8 : _zz_targets_0_bestRequest_id_11);
  assign _zz_targets_0_bestRequest_id_54 = ((! _zz_targets_0_bestRequest_id_17) || (_zz_targets_0_bestRequest_id_14 && (_zz_targets_0_bestRequest_id_16 <= _zz_targets_0_bestRequest_id_13)));
  assign _zz_targets_0_bestRequest_id_55 = (_zz_targets_0_bestRequest_id_54 ? _zz_targets_0_bestRequest_id_13 : _zz_targets_0_bestRequest_id_16);
  assign _zz_targets_0_bestRequest_id_56 = (_zz_targets_0_bestRequest_id_54 ? _zz_targets_0_bestRequest_id_14 : _zz_targets_0_bestRequest_id_17);
  assign _zz_targets_0_bestRequest_id_57 = ((! _zz_targets_0_bestRequest_id_23) || (_zz_targets_0_bestRequest_id_20 && (_zz_targets_0_bestRequest_id_22 <= _zz_targets_0_bestRequest_id_19)));
  assign _zz_targets_0_bestRequest_id_58 = (_zz_targets_0_bestRequest_id_57 ? _zz_targets_0_bestRequest_id_19 : _zz_targets_0_bestRequest_id_22);
  assign _zz_targets_0_bestRequest_id_59 = (_zz_targets_0_bestRequest_id_57 ? _zz_targets_0_bestRequest_id_20 : _zz_targets_0_bestRequest_id_23);
  assign _zz_targets_0_bestRequest_id_60 = ((! _zz_targets_0_bestRequest_id_29) || (_zz_targets_0_bestRequest_id_26 && (_zz_targets_0_bestRequest_id_28 <= _zz_targets_0_bestRequest_id_25)));
  assign _zz_targets_0_bestRequest_id_61 = (_zz_targets_0_bestRequest_id_60 ? _zz_targets_0_bestRequest_id_25 : _zz_targets_0_bestRequest_id_28);
  assign _zz_targets_0_bestRequest_id_62 = (_zz_targets_0_bestRequest_id_60 ? _zz_targets_0_bestRequest_id_26 : _zz_targets_0_bestRequest_id_29);
  assign _zz_targets_0_bestRequest_id_63 = ((! _zz_targets_0_bestRequest_id_35) || (_zz_targets_0_bestRequest_id_32 && (_zz_targets_0_bestRequest_id_34 <= _zz_targets_0_bestRequest_id_31)));
  assign _zz_targets_0_bestRequest_id_64 = (_zz_targets_0_bestRequest_id_63 ? _zz_targets_0_bestRequest_id_31 : _zz_targets_0_bestRequest_id_34);
  assign _zz_targets_0_bestRequest_id_65 = (_zz_targets_0_bestRequest_id_63 ? _zz_targets_0_bestRequest_id_32 : _zz_targets_0_bestRequest_id_35);
  assign _zz_targets_0_bestRequest_id_66 = ((! _zz_targets_0_bestRequest_id_41) || (_zz_targets_0_bestRequest_id_38 && (_zz_targets_0_bestRequest_id_40 <= _zz_targets_0_bestRequest_id_37)));
  assign _zz_targets_0_bestRequest_id_67 = (_zz_targets_0_bestRequest_id_66 ? _zz_targets_0_bestRequest_id_37 : _zz_targets_0_bestRequest_id_40);
  assign _zz_targets_0_bestRequest_id_68 = (_zz_targets_0_bestRequest_id_66 ? _zz_targets_0_bestRequest_id_38 : _zz_targets_0_bestRequest_id_41);
  assign _zz_targets_0_bestRequest_id_69 = ((! _zz_targets_0_bestRequest_id_47) || (_zz_targets_0_bestRequest_id_44 && (_zz_targets_0_bestRequest_id_46 <= _zz_targets_0_bestRequest_id_43)));
  assign _zz_targets_0_bestRequest_id_70 = (_zz_targets_0_bestRequest_id_69 ? _zz_targets_0_bestRequest_id_43 : _zz_targets_0_bestRequest_id_46);
  assign _zz_targets_0_bestRequest_id_71 = (_zz_targets_0_bestRequest_id_69 ? _zz_targets_0_bestRequest_id_44 : _zz_targets_0_bestRequest_id_47);
  assign _zz_targets_0_bestRequest_id_72 = ((! _zz_targets_0_bestRequest_id_53) || (_zz_targets_0_bestRequest_id_50 && (_zz_targets_0_bestRequest_id_52 <= _zz_targets_0_bestRequest_id_49)));
  assign _zz_targets_0_bestRequest_priority = (_zz_targets_0_bestRequest_id_72 ? _zz_targets_0_bestRequest_id_49 : _zz_targets_0_bestRequest_id_52);
  assign _zz_targets_0_bestRequest_id_73 = (_zz_targets_0_bestRequest_id_72 ? _zz_targets_0_bestRequest_id_50 : _zz_targets_0_bestRequest_id_53);
  assign _zz_targets_0_bestRequest_id_74 = ((! _zz_targets_0_bestRequest_id_59) || (_zz_targets_0_bestRequest_id_56 && (_zz_targets_0_bestRequest_id_58 <= _zz_targets_0_bestRequest_id_55)));
  assign _zz_targets_0_bestRequest_priority_1 = (_zz_targets_0_bestRequest_id_74 ? _zz_targets_0_bestRequest_id_55 : _zz_targets_0_bestRequest_id_58);
  assign _zz_targets_0_bestRequest_id_75 = (_zz_targets_0_bestRequest_id_74 ? _zz_targets_0_bestRequest_id_56 : _zz_targets_0_bestRequest_id_59);
  assign _zz_targets_0_bestRequest_id_76 = ((! _zz_targets_0_bestRequest_id_65) || (_zz_targets_0_bestRequest_id_62 && (_zz_targets_0_bestRequest_id_64 <= _zz_targets_0_bestRequest_id_61)));
  assign _zz_targets_0_bestRequest_priority_2 = (_zz_targets_0_bestRequest_id_76 ? _zz_targets_0_bestRequest_id_61 : _zz_targets_0_bestRequest_id_64);
  assign _zz_targets_0_bestRequest_id_77 = (_zz_targets_0_bestRequest_id_76 ? _zz_targets_0_bestRequest_id_62 : _zz_targets_0_bestRequest_id_65);
  assign _zz_targets_0_bestRequest_id_78 = ((! _zz_targets_0_bestRequest_id_71) || (_zz_targets_0_bestRequest_id_68 && (_zz_targets_0_bestRequest_id_70 <= _zz_targets_0_bestRequest_id_67)));
  assign _zz_targets_0_bestRequest_priority_3 = (_zz_targets_0_bestRequest_id_78 ? _zz_targets_0_bestRequest_id_67 : _zz_targets_0_bestRequest_id_70);
  assign _zz_targets_0_bestRequest_id_79 = (_zz_targets_0_bestRequest_id_78 ? _zz_targets_0_bestRequest_id_68 : _zz_targets_0_bestRequest_id_71);
  assign _zz_targets_0_bestRequest_id_80 = ((! _zz_targets_0_bestRequest_id_75) || (_zz_targets_0_bestRequest_id_73 && (_zz_targets_0_bestRequest_priority_1 <= _zz_targets_0_bestRequest_priority)));
  assign _zz_targets_0_bestRequest_priority_4 = (_zz_targets_0_bestRequest_id_80 ? _zz_targets_0_bestRequest_priority : _zz_targets_0_bestRequest_priority_1);
  assign _zz_targets_0_bestRequest_valid = (_zz_targets_0_bestRequest_id_80 ? _zz_targets_0_bestRequest_id_73 : _zz_targets_0_bestRequest_id_75);
  assign _zz_targets_0_bestRequest_id_81 = ((! _zz_targets_0_bestRequest_id_79) || (_zz_targets_0_bestRequest_id_77 && (_zz_targets_0_bestRequest_priority_3 <= _zz_targets_0_bestRequest_priority_2)));
  assign _zz_targets_0_bestRequest_priority_5 = (_zz_targets_0_bestRequest_id_81 ? _zz_targets_0_bestRequest_priority_2 : _zz_targets_0_bestRequest_priority_3);
  assign _zz_targets_0_bestRequest_valid_1 = (_zz_targets_0_bestRequest_id_81 ? _zz_targets_0_bestRequest_id_77 : _zz_targets_0_bestRequest_id_79);
  assign _zz_targets_0_bestRequest_priority_6 = ((! _zz_targets_0_bestRequest_valid_1) || (_zz_targets_0_bestRequest_valid && (_zz_targets_0_bestRequest_priority_5 <= _zz_targets_0_bestRequest_priority_4)));
  assign targets_0_iep = (targets_0_threshold < targets_0_bestRequest_priority);
  assign targets_0_claim = (targets_0_iep ? targets_0_bestRequest_id : 5'h0);
  assign targets_1_requests_0_priority = 2'b00;
  assign targets_1_requests_0_id = 5'h0;
  assign targets_1_requests_0_valid = 1'b1;
  assign targets_1_requests_1_priority = gateways_0_priority;
  assign targets_1_requests_1_id = 5'h01;
  assign targets_1_requests_1_valid = (gateways_0_ip && targets_1_ie_0);
  assign targets_1_requests_2_priority = gateways_1_priority;
  assign targets_1_requests_2_id = 5'h02;
  assign targets_1_requests_2_valid = (gateways_1_ip && targets_1_ie_1);
  assign targets_1_requests_3_priority = gateways_2_priority;
  assign targets_1_requests_3_id = 5'h03;
  assign targets_1_requests_3_valid = (gateways_2_ip && targets_1_ie_2);
  assign targets_1_requests_4_priority = gateways_3_priority;
  assign targets_1_requests_4_id = 5'h04;
  assign targets_1_requests_4_valid = (gateways_3_ip && targets_1_ie_3);
  assign targets_1_requests_5_priority = gateways_4_priority;
  assign targets_1_requests_5_id = 5'h05;
  assign targets_1_requests_5_valid = (gateways_4_ip && targets_1_ie_4);
  assign targets_1_requests_6_priority = gateways_5_priority;
  assign targets_1_requests_6_id = 5'h06;
  assign targets_1_requests_6_valid = (gateways_5_ip && targets_1_ie_5);
  assign targets_1_requests_7_priority = gateways_6_priority;
  assign targets_1_requests_7_id = 5'h07;
  assign targets_1_requests_7_valid = (gateways_6_ip && targets_1_ie_6);
  assign targets_1_requests_8_priority = gateways_7_priority;
  assign targets_1_requests_8_id = 5'h08;
  assign targets_1_requests_8_valid = (gateways_7_ip && targets_1_ie_7);
  assign targets_1_requests_9_priority = gateways_8_priority;
  assign targets_1_requests_9_id = 5'h09;
  assign targets_1_requests_9_valid = (gateways_8_ip && targets_1_ie_8);
  assign targets_1_requests_10_priority = gateways_9_priority;
  assign targets_1_requests_10_id = 5'h0a;
  assign targets_1_requests_10_valid = (gateways_9_ip && targets_1_ie_9);
  assign targets_1_requests_11_priority = gateways_10_priority;
  assign targets_1_requests_11_id = 5'h0b;
  assign targets_1_requests_11_valid = (gateways_10_ip && targets_1_ie_10);
  assign targets_1_requests_12_priority = gateways_11_priority;
  assign targets_1_requests_12_id = 5'h0c;
  assign targets_1_requests_12_valid = (gateways_11_ip && targets_1_ie_11);
  assign targets_1_requests_13_priority = gateways_12_priority;
  assign targets_1_requests_13_id = 5'h0d;
  assign targets_1_requests_13_valid = (gateways_12_ip && targets_1_ie_12);
  assign targets_1_requests_14_priority = gateways_13_priority;
  assign targets_1_requests_14_id = 5'h0e;
  assign targets_1_requests_14_valid = (gateways_13_ip && targets_1_ie_13);
  assign targets_1_requests_15_priority = gateways_14_priority;
  assign targets_1_requests_15_id = 5'h0f;
  assign targets_1_requests_15_valid = (gateways_14_ip && targets_1_ie_14);
  assign targets_1_requests_16_priority = gateways_15_priority;
  assign targets_1_requests_16_id = 5'h10;
  assign targets_1_requests_16_valid = (gateways_15_ip && targets_1_ie_15);
  assign targets_1_requests_17_priority = gateways_16_priority;
  assign targets_1_requests_17_id = 5'h11;
  assign targets_1_requests_17_valid = (gateways_16_ip && targets_1_ie_16);
  assign targets_1_requests_18_priority = gateways_17_priority;
  assign targets_1_requests_18_id = 5'h12;
  assign targets_1_requests_18_valid = (gateways_17_ip && targets_1_ie_17);
  assign targets_1_requests_19_priority = gateways_18_priority;
  assign targets_1_requests_19_id = 5'h13;
  assign targets_1_requests_19_valid = (gateways_18_ip && targets_1_ie_18);
  assign targets_1_requests_20_priority = gateways_19_priority;
  assign targets_1_requests_20_id = 5'h14;
  assign targets_1_requests_20_valid = (gateways_19_ip && targets_1_ie_19);
  assign targets_1_requests_21_priority = gateways_20_priority;
  assign targets_1_requests_21_id = 5'h15;
  assign targets_1_requests_21_valid = (gateways_20_ip && targets_1_ie_20);
  assign targets_1_requests_22_priority = gateways_21_priority;
  assign targets_1_requests_22_id = 5'h16;
  assign targets_1_requests_22_valid = (gateways_21_ip && targets_1_ie_21);
  assign targets_1_requests_23_priority = gateways_22_priority;
  assign targets_1_requests_23_id = 5'h17;
  assign targets_1_requests_23_valid = (gateways_22_ip && targets_1_ie_22);
  assign targets_1_requests_24_priority = gateways_23_priority;
  assign targets_1_requests_24_id = 5'h18;
  assign targets_1_requests_24_valid = (gateways_23_ip && targets_1_ie_23);
  assign targets_1_requests_25_priority = gateways_24_priority;
  assign targets_1_requests_25_id = 5'h19;
  assign targets_1_requests_25_valid = (gateways_24_ip && targets_1_ie_24);
  assign targets_1_requests_26_priority = gateways_25_priority;
  assign targets_1_requests_26_id = 5'h1a;
  assign targets_1_requests_26_valid = (gateways_25_ip && targets_1_ie_25);
  assign targets_1_requests_27_priority = gateways_26_priority;
  assign targets_1_requests_27_id = 5'h1b;
  assign targets_1_requests_27_valid = (gateways_26_ip && targets_1_ie_26);
  assign targets_1_requests_28_priority = gateways_27_priority;
  assign targets_1_requests_28_id = 5'h1c;
  assign targets_1_requests_28_valid = (gateways_27_ip && targets_1_ie_27);
  assign targets_1_requests_29_priority = gateways_28_priority;
  assign targets_1_requests_29_id = 5'h1d;
  assign targets_1_requests_29_valid = (gateways_28_ip && targets_1_ie_28);
  assign targets_1_requests_30_priority = gateways_29_priority;
  assign targets_1_requests_30_id = 5'h1e;
  assign targets_1_requests_30_valid = (gateways_29_ip && targets_1_ie_29);
  assign targets_1_requests_31_priority = gateways_30_priority;
  assign targets_1_requests_31_id = 5'h1f;
  assign targets_1_requests_31_valid = (gateways_30_ip && targets_1_ie_30);
  assign _zz_targets_1_bestRequest_id = ((! targets_1_requests_1_valid) || (targets_1_requests_0_valid && (targets_1_requests_1_priority <= targets_1_requests_0_priority)));
  assign _zz_targets_1_bestRequest_id_1 = (_zz_targets_1_bestRequest_id ? targets_1_requests_0_priority : targets_1_requests_1_priority);
  assign _zz_targets_1_bestRequest_id_2 = (_zz_targets_1_bestRequest_id ? targets_1_requests_0_valid : targets_1_requests_1_valid);
  assign _zz_targets_1_bestRequest_id_3 = ((! targets_1_requests_3_valid) || (targets_1_requests_2_valid && (targets_1_requests_3_priority <= targets_1_requests_2_priority)));
  assign _zz_targets_1_bestRequest_id_4 = (_zz_targets_1_bestRequest_id_3 ? targets_1_requests_2_priority : targets_1_requests_3_priority);
  assign _zz_targets_1_bestRequest_id_5 = (_zz_targets_1_bestRequest_id_3 ? targets_1_requests_2_valid : targets_1_requests_3_valid);
  assign _zz_targets_1_bestRequest_id_6 = ((! targets_1_requests_5_valid) || (targets_1_requests_4_valid && (targets_1_requests_5_priority <= targets_1_requests_4_priority)));
  assign _zz_targets_1_bestRequest_id_7 = (_zz_targets_1_bestRequest_id_6 ? targets_1_requests_4_priority : targets_1_requests_5_priority);
  assign _zz_targets_1_bestRequest_id_8 = (_zz_targets_1_bestRequest_id_6 ? targets_1_requests_4_valid : targets_1_requests_5_valid);
  assign _zz_targets_1_bestRequest_id_9 = ((! targets_1_requests_7_valid) || (targets_1_requests_6_valid && (targets_1_requests_7_priority <= targets_1_requests_6_priority)));
  assign _zz_targets_1_bestRequest_id_10 = (_zz_targets_1_bestRequest_id_9 ? targets_1_requests_6_priority : targets_1_requests_7_priority);
  assign _zz_targets_1_bestRequest_id_11 = (_zz_targets_1_bestRequest_id_9 ? targets_1_requests_6_valid : targets_1_requests_7_valid);
  assign _zz_targets_1_bestRequest_id_12 = ((! targets_1_requests_9_valid) || (targets_1_requests_8_valid && (targets_1_requests_9_priority <= targets_1_requests_8_priority)));
  assign _zz_targets_1_bestRequest_id_13 = (_zz_targets_1_bestRequest_id_12 ? targets_1_requests_8_priority : targets_1_requests_9_priority);
  assign _zz_targets_1_bestRequest_id_14 = (_zz_targets_1_bestRequest_id_12 ? targets_1_requests_8_valid : targets_1_requests_9_valid);
  assign _zz_targets_1_bestRequest_id_15 = ((! targets_1_requests_11_valid) || (targets_1_requests_10_valid && (targets_1_requests_11_priority <= targets_1_requests_10_priority)));
  assign _zz_targets_1_bestRequest_id_16 = (_zz_targets_1_bestRequest_id_15 ? targets_1_requests_10_priority : targets_1_requests_11_priority);
  assign _zz_targets_1_bestRequest_id_17 = (_zz_targets_1_bestRequest_id_15 ? targets_1_requests_10_valid : targets_1_requests_11_valid);
  assign _zz_targets_1_bestRequest_id_18 = ((! targets_1_requests_13_valid) || (targets_1_requests_12_valid && (targets_1_requests_13_priority <= targets_1_requests_12_priority)));
  assign _zz_targets_1_bestRequest_id_19 = (_zz_targets_1_bestRequest_id_18 ? targets_1_requests_12_priority : targets_1_requests_13_priority);
  assign _zz_targets_1_bestRequest_id_20 = (_zz_targets_1_bestRequest_id_18 ? targets_1_requests_12_valid : targets_1_requests_13_valid);
  assign _zz_targets_1_bestRequest_id_21 = ((! targets_1_requests_15_valid) || (targets_1_requests_14_valid && (targets_1_requests_15_priority <= targets_1_requests_14_priority)));
  assign _zz_targets_1_bestRequest_id_22 = (_zz_targets_1_bestRequest_id_21 ? targets_1_requests_14_priority : targets_1_requests_15_priority);
  assign _zz_targets_1_bestRequest_id_23 = (_zz_targets_1_bestRequest_id_21 ? targets_1_requests_14_valid : targets_1_requests_15_valid);
  assign _zz_targets_1_bestRequest_id_24 = ((! targets_1_requests_17_valid) || (targets_1_requests_16_valid && (targets_1_requests_17_priority <= targets_1_requests_16_priority)));
  assign _zz_targets_1_bestRequest_id_25 = (_zz_targets_1_bestRequest_id_24 ? targets_1_requests_16_priority : targets_1_requests_17_priority);
  assign _zz_targets_1_bestRequest_id_26 = (_zz_targets_1_bestRequest_id_24 ? targets_1_requests_16_valid : targets_1_requests_17_valid);
  assign _zz_targets_1_bestRequest_id_27 = ((! targets_1_requests_19_valid) || (targets_1_requests_18_valid && (targets_1_requests_19_priority <= targets_1_requests_18_priority)));
  assign _zz_targets_1_bestRequest_id_28 = (_zz_targets_1_bestRequest_id_27 ? targets_1_requests_18_priority : targets_1_requests_19_priority);
  assign _zz_targets_1_bestRequest_id_29 = (_zz_targets_1_bestRequest_id_27 ? targets_1_requests_18_valid : targets_1_requests_19_valid);
  assign _zz_targets_1_bestRequest_id_30 = ((! targets_1_requests_21_valid) || (targets_1_requests_20_valid && (targets_1_requests_21_priority <= targets_1_requests_20_priority)));
  assign _zz_targets_1_bestRequest_id_31 = (_zz_targets_1_bestRequest_id_30 ? targets_1_requests_20_priority : targets_1_requests_21_priority);
  assign _zz_targets_1_bestRequest_id_32 = (_zz_targets_1_bestRequest_id_30 ? targets_1_requests_20_valid : targets_1_requests_21_valid);
  assign _zz_targets_1_bestRequest_id_33 = ((! targets_1_requests_23_valid) || (targets_1_requests_22_valid && (targets_1_requests_23_priority <= targets_1_requests_22_priority)));
  assign _zz_targets_1_bestRequest_id_34 = (_zz_targets_1_bestRequest_id_33 ? targets_1_requests_22_priority : targets_1_requests_23_priority);
  assign _zz_targets_1_bestRequest_id_35 = (_zz_targets_1_bestRequest_id_33 ? targets_1_requests_22_valid : targets_1_requests_23_valid);
  assign _zz_targets_1_bestRequest_id_36 = ((! targets_1_requests_25_valid) || (targets_1_requests_24_valid && (targets_1_requests_25_priority <= targets_1_requests_24_priority)));
  assign _zz_targets_1_bestRequest_id_37 = (_zz_targets_1_bestRequest_id_36 ? targets_1_requests_24_priority : targets_1_requests_25_priority);
  assign _zz_targets_1_bestRequest_id_38 = (_zz_targets_1_bestRequest_id_36 ? targets_1_requests_24_valid : targets_1_requests_25_valid);
  assign _zz_targets_1_bestRequest_id_39 = ((! targets_1_requests_27_valid) || (targets_1_requests_26_valid && (targets_1_requests_27_priority <= targets_1_requests_26_priority)));
  assign _zz_targets_1_bestRequest_id_40 = (_zz_targets_1_bestRequest_id_39 ? targets_1_requests_26_priority : targets_1_requests_27_priority);
  assign _zz_targets_1_bestRequest_id_41 = (_zz_targets_1_bestRequest_id_39 ? targets_1_requests_26_valid : targets_1_requests_27_valid);
  assign _zz_targets_1_bestRequest_id_42 = ((! targets_1_requests_29_valid) || (targets_1_requests_28_valid && (targets_1_requests_29_priority <= targets_1_requests_28_priority)));
  assign _zz_targets_1_bestRequest_id_43 = (_zz_targets_1_bestRequest_id_42 ? targets_1_requests_28_priority : targets_1_requests_29_priority);
  assign _zz_targets_1_bestRequest_id_44 = (_zz_targets_1_bestRequest_id_42 ? targets_1_requests_28_valid : targets_1_requests_29_valid);
  assign _zz_targets_1_bestRequest_id_45 = ((! targets_1_requests_31_valid) || (targets_1_requests_30_valid && (targets_1_requests_31_priority <= targets_1_requests_30_priority)));
  assign _zz_targets_1_bestRequest_id_46 = (_zz_targets_1_bestRequest_id_45 ? targets_1_requests_30_priority : targets_1_requests_31_priority);
  assign _zz_targets_1_bestRequest_id_47 = (_zz_targets_1_bestRequest_id_45 ? targets_1_requests_30_valid : targets_1_requests_31_valid);
  assign _zz_targets_1_bestRequest_id_48 = ((! _zz_targets_1_bestRequest_id_5) || (_zz_targets_1_bestRequest_id_2 && (_zz_targets_1_bestRequest_id_4 <= _zz_targets_1_bestRequest_id_1)));
  assign _zz_targets_1_bestRequest_id_49 = (_zz_targets_1_bestRequest_id_48 ? _zz_targets_1_bestRequest_id_1 : _zz_targets_1_bestRequest_id_4);
  assign _zz_targets_1_bestRequest_id_50 = (_zz_targets_1_bestRequest_id_48 ? _zz_targets_1_bestRequest_id_2 : _zz_targets_1_bestRequest_id_5);
  assign _zz_targets_1_bestRequest_id_51 = ((! _zz_targets_1_bestRequest_id_11) || (_zz_targets_1_bestRequest_id_8 && (_zz_targets_1_bestRequest_id_10 <= _zz_targets_1_bestRequest_id_7)));
  assign _zz_targets_1_bestRequest_id_52 = (_zz_targets_1_bestRequest_id_51 ? _zz_targets_1_bestRequest_id_7 : _zz_targets_1_bestRequest_id_10);
  assign _zz_targets_1_bestRequest_id_53 = (_zz_targets_1_bestRequest_id_51 ? _zz_targets_1_bestRequest_id_8 : _zz_targets_1_bestRequest_id_11);
  assign _zz_targets_1_bestRequest_id_54 = ((! _zz_targets_1_bestRequest_id_17) || (_zz_targets_1_bestRequest_id_14 && (_zz_targets_1_bestRequest_id_16 <= _zz_targets_1_bestRequest_id_13)));
  assign _zz_targets_1_bestRequest_id_55 = (_zz_targets_1_bestRequest_id_54 ? _zz_targets_1_bestRequest_id_13 : _zz_targets_1_bestRequest_id_16);
  assign _zz_targets_1_bestRequest_id_56 = (_zz_targets_1_bestRequest_id_54 ? _zz_targets_1_bestRequest_id_14 : _zz_targets_1_bestRequest_id_17);
  assign _zz_targets_1_bestRequest_id_57 = ((! _zz_targets_1_bestRequest_id_23) || (_zz_targets_1_bestRequest_id_20 && (_zz_targets_1_bestRequest_id_22 <= _zz_targets_1_bestRequest_id_19)));
  assign _zz_targets_1_bestRequest_id_58 = (_zz_targets_1_bestRequest_id_57 ? _zz_targets_1_bestRequest_id_19 : _zz_targets_1_bestRequest_id_22);
  assign _zz_targets_1_bestRequest_id_59 = (_zz_targets_1_bestRequest_id_57 ? _zz_targets_1_bestRequest_id_20 : _zz_targets_1_bestRequest_id_23);
  assign _zz_targets_1_bestRequest_id_60 = ((! _zz_targets_1_bestRequest_id_29) || (_zz_targets_1_bestRequest_id_26 && (_zz_targets_1_bestRequest_id_28 <= _zz_targets_1_bestRequest_id_25)));
  assign _zz_targets_1_bestRequest_id_61 = (_zz_targets_1_bestRequest_id_60 ? _zz_targets_1_bestRequest_id_25 : _zz_targets_1_bestRequest_id_28);
  assign _zz_targets_1_bestRequest_id_62 = (_zz_targets_1_bestRequest_id_60 ? _zz_targets_1_bestRequest_id_26 : _zz_targets_1_bestRequest_id_29);
  assign _zz_targets_1_bestRequest_id_63 = ((! _zz_targets_1_bestRequest_id_35) || (_zz_targets_1_bestRequest_id_32 && (_zz_targets_1_bestRequest_id_34 <= _zz_targets_1_bestRequest_id_31)));
  assign _zz_targets_1_bestRequest_id_64 = (_zz_targets_1_bestRequest_id_63 ? _zz_targets_1_bestRequest_id_31 : _zz_targets_1_bestRequest_id_34);
  assign _zz_targets_1_bestRequest_id_65 = (_zz_targets_1_bestRequest_id_63 ? _zz_targets_1_bestRequest_id_32 : _zz_targets_1_bestRequest_id_35);
  assign _zz_targets_1_bestRequest_id_66 = ((! _zz_targets_1_bestRequest_id_41) || (_zz_targets_1_bestRequest_id_38 && (_zz_targets_1_bestRequest_id_40 <= _zz_targets_1_bestRequest_id_37)));
  assign _zz_targets_1_bestRequest_id_67 = (_zz_targets_1_bestRequest_id_66 ? _zz_targets_1_bestRequest_id_37 : _zz_targets_1_bestRequest_id_40);
  assign _zz_targets_1_bestRequest_id_68 = (_zz_targets_1_bestRequest_id_66 ? _zz_targets_1_bestRequest_id_38 : _zz_targets_1_bestRequest_id_41);
  assign _zz_targets_1_bestRequest_id_69 = ((! _zz_targets_1_bestRequest_id_47) || (_zz_targets_1_bestRequest_id_44 && (_zz_targets_1_bestRequest_id_46 <= _zz_targets_1_bestRequest_id_43)));
  assign _zz_targets_1_bestRequest_id_70 = (_zz_targets_1_bestRequest_id_69 ? _zz_targets_1_bestRequest_id_43 : _zz_targets_1_bestRequest_id_46);
  assign _zz_targets_1_bestRequest_id_71 = (_zz_targets_1_bestRequest_id_69 ? _zz_targets_1_bestRequest_id_44 : _zz_targets_1_bestRequest_id_47);
  assign _zz_targets_1_bestRequest_id_72 = ((! _zz_targets_1_bestRequest_id_53) || (_zz_targets_1_bestRequest_id_50 && (_zz_targets_1_bestRequest_id_52 <= _zz_targets_1_bestRequest_id_49)));
  assign _zz_targets_1_bestRequest_priority = (_zz_targets_1_bestRequest_id_72 ? _zz_targets_1_bestRequest_id_49 : _zz_targets_1_bestRequest_id_52);
  assign _zz_targets_1_bestRequest_id_73 = (_zz_targets_1_bestRequest_id_72 ? _zz_targets_1_bestRequest_id_50 : _zz_targets_1_bestRequest_id_53);
  assign _zz_targets_1_bestRequest_id_74 = ((! _zz_targets_1_bestRequest_id_59) || (_zz_targets_1_bestRequest_id_56 && (_zz_targets_1_bestRequest_id_58 <= _zz_targets_1_bestRequest_id_55)));
  assign _zz_targets_1_bestRequest_priority_1 = (_zz_targets_1_bestRequest_id_74 ? _zz_targets_1_bestRequest_id_55 : _zz_targets_1_bestRequest_id_58);
  assign _zz_targets_1_bestRequest_id_75 = (_zz_targets_1_bestRequest_id_74 ? _zz_targets_1_bestRequest_id_56 : _zz_targets_1_bestRequest_id_59);
  assign _zz_targets_1_bestRequest_id_76 = ((! _zz_targets_1_bestRequest_id_65) || (_zz_targets_1_bestRequest_id_62 && (_zz_targets_1_bestRequest_id_64 <= _zz_targets_1_bestRequest_id_61)));
  assign _zz_targets_1_bestRequest_priority_2 = (_zz_targets_1_bestRequest_id_76 ? _zz_targets_1_bestRequest_id_61 : _zz_targets_1_bestRequest_id_64);
  assign _zz_targets_1_bestRequest_id_77 = (_zz_targets_1_bestRequest_id_76 ? _zz_targets_1_bestRequest_id_62 : _zz_targets_1_bestRequest_id_65);
  assign _zz_targets_1_bestRequest_id_78 = ((! _zz_targets_1_bestRequest_id_71) || (_zz_targets_1_bestRequest_id_68 && (_zz_targets_1_bestRequest_id_70 <= _zz_targets_1_bestRequest_id_67)));
  assign _zz_targets_1_bestRequest_priority_3 = (_zz_targets_1_bestRequest_id_78 ? _zz_targets_1_bestRequest_id_67 : _zz_targets_1_bestRequest_id_70);
  assign _zz_targets_1_bestRequest_id_79 = (_zz_targets_1_bestRequest_id_78 ? _zz_targets_1_bestRequest_id_68 : _zz_targets_1_bestRequest_id_71);
  assign _zz_targets_1_bestRequest_id_80 = ((! _zz_targets_1_bestRequest_id_75) || (_zz_targets_1_bestRequest_id_73 && (_zz_targets_1_bestRequest_priority_1 <= _zz_targets_1_bestRequest_priority)));
  assign _zz_targets_1_bestRequest_priority_4 = (_zz_targets_1_bestRequest_id_80 ? _zz_targets_1_bestRequest_priority : _zz_targets_1_bestRequest_priority_1);
  assign _zz_targets_1_bestRequest_valid = (_zz_targets_1_bestRequest_id_80 ? _zz_targets_1_bestRequest_id_73 : _zz_targets_1_bestRequest_id_75);
  assign _zz_targets_1_bestRequest_id_81 = ((! _zz_targets_1_bestRequest_id_79) || (_zz_targets_1_bestRequest_id_77 && (_zz_targets_1_bestRequest_priority_3 <= _zz_targets_1_bestRequest_priority_2)));
  assign _zz_targets_1_bestRequest_priority_5 = (_zz_targets_1_bestRequest_id_81 ? _zz_targets_1_bestRequest_priority_2 : _zz_targets_1_bestRequest_priority_3);
  assign _zz_targets_1_bestRequest_valid_1 = (_zz_targets_1_bestRequest_id_81 ? _zz_targets_1_bestRequest_id_77 : _zz_targets_1_bestRequest_id_79);
  assign _zz_targets_1_bestRequest_priority_6 = ((! _zz_targets_1_bestRequest_valid_1) || (_zz_targets_1_bestRequest_valid && (_zz_targets_1_bestRequest_priority_5 <= _zz_targets_1_bestRequest_priority_4)));
  assign targets_1_iep = (targets_1_threshold < targets_1_bestRequest_priority);
  assign targets_1_claim = (targets_1_iep ? targets_1_bestRequest_id : 5'h0);
  assign io_targets = {targets_1_iep,targets_0_iep};
  assign factory_readErrorFlag = 1'b0;
  assign factory_writeErrorFlag = 1'b0;
  assign factory_askWrite = (io_bus_a_valid && (|{(io_bus_a_payload_opcode == A_PUT_PARTIAL_DATA),(io_bus_a_payload_opcode == A_PUT_FULL_DATA)}));
  assign factory_askRead = (io_bus_a_valid && (|(io_bus_a_payload_opcode == A_GET)));
  assign factory_doWrite = (factory_askWrite && io_bus_a_ready);
  assign factory_doRead = (factory_askRead && io_bus_a_ready);
  assign factory_address = ({2'd0,_zz_factory_address} <<< 2'd2);
  always @(*) begin
    factory_halt = 1'b0;
    if(when_PlicMapper_l122) begin
      factory_halt = 1'b1;
    end
  end

  assign gateways_0_priority = gateways_0_priority_driver;
  assign gateways_1_priority = gateways_1_priority_driver;
  assign gateways_2_priority = gateways_2_priority_driver;
  assign gateways_3_priority = gateways_3_priority_driver;
  assign gateways_4_priority = gateways_4_priority_driver;
  assign gateways_5_priority = gateways_5_priority_driver;
  assign gateways_6_priority = gateways_6_priority_driver;
  assign gateways_7_priority = gateways_7_priority_driver;
  assign gateways_8_priority = gateways_8_priority_driver;
  assign gateways_9_priority = gateways_9_priority_driver;
  assign gateways_10_priority = gateways_10_priority_driver;
  assign gateways_11_priority = gateways_11_priority_driver;
  assign gateways_12_priority = gateways_12_priority_driver;
  assign gateways_13_priority = gateways_13_priority_driver;
  assign gateways_14_priority = gateways_14_priority_driver;
  assign gateways_15_priority = gateways_15_priority_driver;
  assign gateways_16_priority = gateways_16_priority_driver;
  assign gateways_17_priority = gateways_17_priority_driver;
  assign gateways_18_priority = gateways_18_priority_driver;
  assign gateways_19_priority = gateways_19_priority_driver;
  assign gateways_20_priority = gateways_20_priority_driver;
  assign gateways_21_priority = gateways_21_priority_driver;
  assign gateways_22_priority = gateways_22_priority_driver;
  assign gateways_23_priority = gateways_23_priority_driver;
  assign gateways_24_priority = gateways_24_priority_driver;
  assign gateways_25_priority = gateways_25_priority_driver;
  assign gateways_26_priority = gateways_26_priority_driver;
  assign gateways_27_priority = gateways_27_priority_driver;
  assign gateways_28_priority = gateways_28_priority_driver;
  assign gateways_29_priority = gateways_29_priority_driver;
  assign gateways_30_priority = gateways_30_priority_driver;
  always @(*) begin
    mapping_claim_valid = 1'b0;
    case(factory_address)
      22'h200004 : begin
        if(factory_doRead) begin
          mapping_claim_valid = 1'b1;
        end
      end
      22'h201004 : begin
        if(factory_doRead) begin
          mapping_claim_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mapping_claim_payload = 5'bxxxxx;
    case(factory_address)
      22'h200004 : begin
        if(factory_doRead) begin
          mapping_claim_payload = targets_0_claim;
        end
      end
      22'h201004 : begin
        if(factory_doRead) begin
          mapping_claim_payload = targets_1_claim;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mapping_completion_valid = 1'b0;
    if(mapping_targetMapping_0_targetCompletion_valid) begin
      mapping_completion_valid = 1'b1;
    end
    if(mapping_targetMapping_1_targetCompletion_valid) begin
      mapping_completion_valid = 1'b1;
    end
  end

  always @(*) begin
    mapping_completion_payload = 5'bxxxxx;
    if(mapping_targetMapping_0_targetCompletion_valid) begin
      mapping_completion_payload = mapping_targetMapping_0_targetCompletion_payload;
    end
    if(mapping_targetMapping_1_targetCompletion_valid) begin
      mapping_completion_payload = mapping_targetMapping_1_targetCompletion_payload;
    end
  end

  always @(*) begin
    mapping_coherencyStall_willIncrement = 1'b0;
    if(when_PlicMapper_l122) begin
      mapping_coherencyStall_willIncrement = 1'b1;
    end
    if(when_SlaveFactory_l134) begin
      if(factory_askWrite) begin
        mapping_coherencyStall_willIncrement = 1'b1;
      end
      if(factory_askRead) begin
        mapping_coherencyStall_willIncrement = 1'b1;
      end
    end
  end

  assign mapping_coherencyStall_willClear = 1'b0;
  assign mapping_coherencyStall_willOverflowIfInc = (mapping_coherencyStall_value == 1'b1);
  assign mapping_coherencyStall_willOverflow = (mapping_coherencyStall_willOverflowIfInc && mapping_coherencyStall_willIncrement);
  always @(*) begin
    mapping_coherencyStall_valueNext = (mapping_coherencyStall_value + mapping_coherencyStall_willIncrement);
    if(mapping_coherencyStall_willClear) begin
      mapping_coherencyStall_valueNext = 1'b0;
    end
  end

  assign when_PlicMapper_l122 = (mapping_coherencyStall_value != 1'b0);
  assign targets_0_threshold = targets_0_threshold_driver;
  always @(*) begin
    mapping_targetMapping_0_targetCompletion_valid = 1'b0;
    case(factory_address)
      22'h200004 : begin
        if(factory_doWrite) begin
          mapping_targetMapping_0_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign targets_0_ie_0 = targets_0_ie_0_driver;
  assign targets_0_ie_1 = targets_0_ie_1_driver;
  assign targets_0_ie_2 = targets_0_ie_2_driver;
  assign targets_0_ie_3 = targets_0_ie_3_driver;
  assign targets_0_ie_4 = targets_0_ie_4_driver;
  assign targets_0_ie_5 = targets_0_ie_5_driver;
  assign targets_0_ie_6 = targets_0_ie_6_driver;
  assign targets_0_ie_7 = targets_0_ie_7_driver;
  assign targets_0_ie_8 = targets_0_ie_8_driver;
  assign targets_0_ie_9 = targets_0_ie_9_driver;
  assign targets_0_ie_10 = targets_0_ie_10_driver;
  assign targets_0_ie_11 = targets_0_ie_11_driver;
  assign targets_0_ie_12 = targets_0_ie_12_driver;
  assign targets_0_ie_13 = targets_0_ie_13_driver;
  assign targets_0_ie_14 = targets_0_ie_14_driver;
  assign targets_0_ie_15 = targets_0_ie_15_driver;
  assign targets_0_ie_16 = targets_0_ie_16_driver;
  assign targets_0_ie_17 = targets_0_ie_17_driver;
  assign targets_0_ie_18 = targets_0_ie_18_driver;
  assign targets_0_ie_19 = targets_0_ie_19_driver;
  assign targets_0_ie_20 = targets_0_ie_20_driver;
  assign targets_0_ie_21 = targets_0_ie_21_driver;
  assign targets_0_ie_22 = targets_0_ie_22_driver;
  assign targets_0_ie_23 = targets_0_ie_23_driver;
  assign targets_0_ie_24 = targets_0_ie_24_driver;
  assign targets_0_ie_25 = targets_0_ie_25_driver;
  assign targets_0_ie_26 = targets_0_ie_26_driver;
  assign targets_0_ie_27 = targets_0_ie_27_driver;
  assign targets_0_ie_28 = targets_0_ie_28_driver;
  assign targets_0_ie_29 = targets_0_ie_29_driver;
  assign targets_0_ie_30 = targets_0_ie_30_driver;
  assign targets_1_threshold = targets_1_threshold_driver;
  always @(*) begin
    mapping_targetMapping_1_targetCompletion_valid = 1'b0;
    case(factory_address)
      22'h201004 : begin
        if(factory_doWrite) begin
          mapping_targetMapping_1_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign targets_1_ie_0 = targets_1_ie_0_driver;
  assign targets_1_ie_1 = targets_1_ie_1_driver;
  assign targets_1_ie_2 = targets_1_ie_2_driver;
  assign targets_1_ie_3 = targets_1_ie_3_driver;
  assign targets_1_ie_4 = targets_1_ie_4_driver;
  assign targets_1_ie_5 = targets_1_ie_5_driver;
  assign targets_1_ie_6 = targets_1_ie_6_driver;
  assign targets_1_ie_7 = targets_1_ie_7_driver;
  assign targets_1_ie_8 = targets_1_ie_8_driver;
  assign targets_1_ie_9 = targets_1_ie_9_driver;
  assign targets_1_ie_10 = targets_1_ie_10_driver;
  assign targets_1_ie_11 = targets_1_ie_11_driver;
  assign targets_1_ie_12 = targets_1_ie_12_driver;
  assign targets_1_ie_13 = targets_1_ie_13_driver;
  assign targets_1_ie_14 = targets_1_ie_14_driver;
  assign targets_1_ie_15 = targets_1_ie_15_driver;
  assign targets_1_ie_16 = targets_1_ie_16_driver;
  assign targets_1_ie_17 = targets_1_ie_17_driver;
  assign targets_1_ie_18 = targets_1_ie_18_driver;
  assign targets_1_ie_19 = targets_1_ie_19_driver;
  assign targets_1_ie_20 = targets_1_ie_20_driver;
  assign targets_1_ie_21 = targets_1_ie_21_driver;
  assign targets_1_ie_22 = targets_1_ie_22_driver;
  assign targets_1_ie_23 = targets_1_ie_23_driver;
  assign targets_1_ie_24 = targets_1_ie_24_driver;
  assign targets_1_ie_25 = targets_1_ie_25_driver;
  assign targets_1_ie_26 = targets_1_ie_26_driver;
  assign targets_1_ie_27 = targets_1_ie_27_driver;
  assign targets_1_ie_28 = targets_1_ie_28_driver;
  assign targets_1_ie_29 = targets_1_ie_29_driver;
  assign targets_1_ie_30 = targets_1_ie_30_driver;
  assign mapping_targetMapping_0_targetCompletion_payload = io_bus_a_payload_data[4 : 0];
  assign mapping_targetMapping_1_targetCompletion_payload = io_bus_a_payload_data[4 : 0];
  assign io_bus_a_ready = (factory_rspAsync_ready && (! factory_halt));
  assign factory_rspAsync_valid = ((io_bus_a_valid && (! factory_halt)) && 1'b1);
  always @(*) begin
    factory_rspAsync_payload_data = 32'h0;
    case(factory_address)
      22'h000004 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_0_priority;
      end
      22'h001000 : begin
        factory_rspAsync_payload_data[1 : 1] = gateways_0_ip;
        factory_rspAsync_payload_data[2 : 2] = gateways_1_ip;
        factory_rspAsync_payload_data[3 : 3] = gateways_2_ip;
        factory_rspAsync_payload_data[4 : 4] = gateways_3_ip;
        factory_rspAsync_payload_data[5 : 5] = gateways_4_ip;
        factory_rspAsync_payload_data[6 : 6] = gateways_5_ip;
        factory_rspAsync_payload_data[7 : 7] = gateways_6_ip;
        factory_rspAsync_payload_data[8 : 8] = gateways_7_ip;
        factory_rspAsync_payload_data[9 : 9] = gateways_8_ip;
        factory_rspAsync_payload_data[10 : 10] = gateways_9_ip;
        factory_rspAsync_payload_data[11 : 11] = gateways_10_ip;
        factory_rspAsync_payload_data[12 : 12] = gateways_11_ip;
        factory_rspAsync_payload_data[13 : 13] = gateways_12_ip;
        factory_rspAsync_payload_data[14 : 14] = gateways_13_ip;
        factory_rspAsync_payload_data[15 : 15] = gateways_14_ip;
        factory_rspAsync_payload_data[16 : 16] = gateways_15_ip;
        factory_rspAsync_payload_data[17 : 17] = gateways_16_ip;
        factory_rspAsync_payload_data[18 : 18] = gateways_17_ip;
        factory_rspAsync_payload_data[19 : 19] = gateways_18_ip;
        factory_rspAsync_payload_data[20 : 20] = gateways_19_ip;
        factory_rspAsync_payload_data[21 : 21] = gateways_20_ip;
        factory_rspAsync_payload_data[22 : 22] = gateways_21_ip;
        factory_rspAsync_payload_data[23 : 23] = gateways_22_ip;
        factory_rspAsync_payload_data[24 : 24] = gateways_23_ip;
        factory_rspAsync_payload_data[25 : 25] = gateways_24_ip;
        factory_rspAsync_payload_data[26 : 26] = gateways_25_ip;
        factory_rspAsync_payload_data[27 : 27] = gateways_26_ip;
        factory_rspAsync_payload_data[28 : 28] = gateways_27_ip;
        factory_rspAsync_payload_data[29 : 29] = gateways_28_ip;
        factory_rspAsync_payload_data[30 : 30] = gateways_29_ip;
        factory_rspAsync_payload_data[31 : 31] = gateways_30_ip;
      end
      22'h000008 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_1_priority;
      end
      22'h00000c : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_2_priority;
      end
      22'h000010 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_3_priority;
      end
      22'h000014 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_4_priority;
      end
      22'h000018 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_5_priority;
      end
      22'h00001c : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_6_priority;
      end
      22'h000020 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_7_priority;
      end
      22'h000024 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_8_priority;
      end
      22'h000028 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_9_priority;
      end
      22'h00002c : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_10_priority;
      end
      22'h000030 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_11_priority;
      end
      22'h000034 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_12_priority;
      end
      22'h000038 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_13_priority;
      end
      22'h00003c : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_14_priority;
      end
      22'h000040 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_15_priority;
      end
      22'h000044 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_16_priority;
      end
      22'h000048 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_17_priority;
      end
      22'h00004c : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_18_priority;
      end
      22'h000050 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_19_priority;
      end
      22'h000054 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_20_priority;
      end
      22'h000058 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_21_priority;
      end
      22'h00005c : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_22_priority;
      end
      22'h000060 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_23_priority;
      end
      22'h000064 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_24_priority;
      end
      22'h000068 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_25_priority;
      end
      22'h00006c : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_26_priority;
      end
      22'h000070 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_27_priority;
      end
      22'h000074 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_28_priority;
      end
      22'h000078 : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_29_priority;
      end
      22'h00007c : begin
        factory_rspAsync_payload_data[1 : 0] = gateways_30_priority;
      end
      22'h200000 : begin
        factory_rspAsync_payload_data[1 : 0] = targets_0_threshold;
      end
      22'h200004 : begin
        factory_rspAsync_payload_data[4 : 0] = targets_0_claim;
      end
      22'h002000 : begin
        factory_rspAsync_payload_data[1 : 1] = targets_0_ie_0;
        factory_rspAsync_payload_data[2 : 2] = targets_0_ie_1;
        factory_rspAsync_payload_data[3 : 3] = targets_0_ie_2;
        factory_rspAsync_payload_data[4 : 4] = targets_0_ie_3;
        factory_rspAsync_payload_data[5 : 5] = targets_0_ie_4;
        factory_rspAsync_payload_data[6 : 6] = targets_0_ie_5;
        factory_rspAsync_payload_data[7 : 7] = targets_0_ie_6;
        factory_rspAsync_payload_data[8 : 8] = targets_0_ie_7;
        factory_rspAsync_payload_data[9 : 9] = targets_0_ie_8;
        factory_rspAsync_payload_data[10 : 10] = targets_0_ie_9;
        factory_rspAsync_payload_data[11 : 11] = targets_0_ie_10;
        factory_rspAsync_payload_data[12 : 12] = targets_0_ie_11;
        factory_rspAsync_payload_data[13 : 13] = targets_0_ie_12;
        factory_rspAsync_payload_data[14 : 14] = targets_0_ie_13;
        factory_rspAsync_payload_data[15 : 15] = targets_0_ie_14;
        factory_rspAsync_payload_data[16 : 16] = targets_0_ie_15;
        factory_rspAsync_payload_data[17 : 17] = targets_0_ie_16;
        factory_rspAsync_payload_data[18 : 18] = targets_0_ie_17;
        factory_rspAsync_payload_data[19 : 19] = targets_0_ie_18;
        factory_rspAsync_payload_data[20 : 20] = targets_0_ie_19;
        factory_rspAsync_payload_data[21 : 21] = targets_0_ie_20;
        factory_rspAsync_payload_data[22 : 22] = targets_0_ie_21;
        factory_rspAsync_payload_data[23 : 23] = targets_0_ie_22;
        factory_rspAsync_payload_data[24 : 24] = targets_0_ie_23;
        factory_rspAsync_payload_data[25 : 25] = targets_0_ie_24;
        factory_rspAsync_payload_data[26 : 26] = targets_0_ie_25;
        factory_rspAsync_payload_data[27 : 27] = targets_0_ie_26;
        factory_rspAsync_payload_data[28 : 28] = targets_0_ie_27;
        factory_rspAsync_payload_data[29 : 29] = targets_0_ie_28;
        factory_rspAsync_payload_data[30 : 30] = targets_0_ie_29;
        factory_rspAsync_payload_data[31 : 31] = targets_0_ie_30;
      end
      22'h201000 : begin
        factory_rspAsync_payload_data[1 : 0] = targets_1_threshold;
      end
      22'h201004 : begin
        factory_rspAsync_payload_data[4 : 0] = targets_1_claim;
      end
      22'h002080 : begin
        factory_rspAsync_payload_data[1 : 1] = targets_1_ie_0;
        factory_rspAsync_payload_data[2 : 2] = targets_1_ie_1;
        factory_rspAsync_payload_data[3 : 3] = targets_1_ie_2;
        factory_rspAsync_payload_data[4 : 4] = targets_1_ie_3;
        factory_rspAsync_payload_data[5 : 5] = targets_1_ie_4;
        factory_rspAsync_payload_data[6 : 6] = targets_1_ie_5;
        factory_rspAsync_payload_data[7 : 7] = targets_1_ie_6;
        factory_rspAsync_payload_data[8 : 8] = targets_1_ie_7;
        factory_rspAsync_payload_data[9 : 9] = targets_1_ie_8;
        factory_rspAsync_payload_data[10 : 10] = targets_1_ie_9;
        factory_rspAsync_payload_data[11 : 11] = targets_1_ie_10;
        factory_rspAsync_payload_data[12 : 12] = targets_1_ie_11;
        factory_rspAsync_payload_data[13 : 13] = targets_1_ie_12;
        factory_rspAsync_payload_data[14 : 14] = targets_1_ie_13;
        factory_rspAsync_payload_data[15 : 15] = targets_1_ie_14;
        factory_rspAsync_payload_data[16 : 16] = targets_1_ie_15;
        factory_rspAsync_payload_data[17 : 17] = targets_1_ie_16;
        factory_rspAsync_payload_data[18 : 18] = targets_1_ie_17;
        factory_rspAsync_payload_data[19 : 19] = targets_1_ie_18;
        factory_rspAsync_payload_data[20 : 20] = targets_1_ie_19;
        factory_rspAsync_payload_data[21 : 21] = targets_1_ie_20;
        factory_rspAsync_payload_data[22 : 22] = targets_1_ie_21;
        factory_rspAsync_payload_data[23 : 23] = targets_1_ie_22;
        factory_rspAsync_payload_data[24 : 24] = targets_1_ie_23;
        factory_rspAsync_payload_data[25 : 25] = targets_1_ie_24;
        factory_rspAsync_payload_data[26 : 26] = targets_1_ie_25;
        factory_rspAsync_payload_data[27 : 27] = targets_1_ie_26;
        factory_rspAsync_payload_data[28 : 28] = targets_1_ie_27;
        factory_rspAsync_payload_data[29 : 29] = targets_1_ie_28;
        factory_rspAsync_payload_data[30 : 30] = targets_1_ie_29;
        factory_rspAsync_payload_data[31 : 31] = targets_1_ie_30;
      end
      default : begin
      end
    endcase
  end

  assign _zz_factory_rspAsync_payload_opcode = ((|(io_bus_a_payload_opcode == A_GET)) ? D_ACCESS_ACK_DATA : D_ACCESS_ACK);
  assign factory_rspAsync_payload_opcode = _zz_factory_rspAsync_payload_opcode;
  assign factory_rspAsync_payload_param = 3'b000;
  assign factory_rspAsync_payload_source = io_bus_a_payload_source;
  assign factory_rspAsync_payload_size = io_bus_a_payload_size;
  assign factory_rspAsync_payload_corrupt = 1'b0;
  assign factory_rspAsync_payload_denied = 1'b0;
  always @(*) begin
    factory_rspAsync_ready = factory_rspAsync_stage_ready;
    if(when_Stream_l399) begin
      factory_rspAsync_ready = 1'b1;
    end
  end

  assign when_Stream_l399 = (! factory_rspAsync_stage_valid);
  assign factory_rspAsync_stage_valid = factory_rspAsync_rValid;
  assign factory_rspAsync_stage_payload_opcode = factory_rspAsync_rData_opcode;
  assign factory_rspAsync_stage_payload_param = factory_rspAsync_rData_param;
  assign factory_rspAsync_stage_payload_source = factory_rspAsync_rData_source;
  assign factory_rspAsync_stage_payload_size = factory_rspAsync_rData_size;
  assign factory_rspAsync_stage_payload_denied = factory_rspAsync_rData_denied;
  assign factory_rspAsync_stage_payload_data = factory_rspAsync_rData_data;
  assign factory_rspAsync_stage_payload_corrupt = factory_rspAsync_rData_corrupt;
  assign io_bus_d_valid = factory_rspAsync_stage_valid;
  assign factory_rspAsync_stage_ready = io_bus_d_ready;
  assign io_bus_d_payload_opcode = factory_rspAsync_stage_payload_opcode;
  assign io_bus_d_payload_param = factory_rspAsync_stage_payload_param;
  assign io_bus_d_payload_source = factory_rspAsync_stage_payload_source;
  assign io_bus_d_payload_size = factory_rspAsync_stage_payload_size;
  assign io_bus_d_payload_denied = factory_rspAsync_stage_payload_denied;
  assign io_bus_d_payload_data = factory_rspAsync_stage_payload_data;
  assign io_bus_d_payload_corrupt = factory_rspAsync_stage_payload_corrupt;
  assign when_SlaveFactory_l134 = 1'b1;
  always @(posedge litex_clk or posedge litex_reset) begin
    if(litex_reset) begin
      gateways_0_ip <= 1'b0;
      gateways_0_waitCompletion <= 1'b0;
      gateways_1_ip <= 1'b0;
      gateways_1_waitCompletion <= 1'b0;
      gateways_2_ip <= 1'b0;
      gateways_2_waitCompletion <= 1'b0;
      gateways_3_ip <= 1'b0;
      gateways_3_waitCompletion <= 1'b0;
      gateways_4_ip <= 1'b0;
      gateways_4_waitCompletion <= 1'b0;
      gateways_5_ip <= 1'b0;
      gateways_5_waitCompletion <= 1'b0;
      gateways_6_ip <= 1'b0;
      gateways_6_waitCompletion <= 1'b0;
      gateways_7_ip <= 1'b0;
      gateways_7_waitCompletion <= 1'b0;
      gateways_8_ip <= 1'b0;
      gateways_8_waitCompletion <= 1'b0;
      gateways_9_ip <= 1'b0;
      gateways_9_waitCompletion <= 1'b0;
      gateways_10_ip <= 1'b0;
      gateways_10_waitCompletion <= 1'b0;
      gateways_11_ip <= 1'b0;
      gateways_11_waitCompletion <= 1'b0;
      gateways_12_ip <= 1'b0;
      gateways_12_waitCompletion <= 1'b0;
      gateways_13_ip <= 1'b0;
      gateways_13_waitCompletion <= 1'b0;
      gateways_14_ip <= 1'b0;
      gateways_14_waitCompletion <= 1'b0;
      gateways_15_ip <= 1'b0;
      gateways_15_waitCompletion <= 1'b0;
      gateways_16_ip <= 1'b0;
      gateways_16_waitCompletion <= 1'b0;
      gateways_17_ip <= 1'b0;
      gateways_17_waitCompletion <= 1'b0;
      gateways_18_ip <= 1'b0;
      gateways_18_waitCompletion <= 1'b0;
      gateways_19_ip <= 1'b0;
      gateways_19_waitCompletion <= 1'b0;
      gateways_20_ip <= 1'b0;
      gateways_20_waitCompletion <= 1'b0;
      gateways_21_ip <= 1'b0;
      gateways_21_waitCompletion <= 1'b0;
      gateways_22_ip <= 1'b0;
      gateways_22_waitCompletion <= 1'b0;
      gateways_23_ip <= 1'b0;
      gateways_23_waitCompletion <= 1'b0;
      gateways_24_ip <= 1'b0;
      gateways_24_waitCompletion <= 1'b0;
      gateways_25_ip <= 1'b0;
      gateways_25_waitCompletion <= 1'b0;
      gateways_26_ip <= 1'b0;
      gateways_26_waitCompletion <= 1'b0;
      gateways_27_ip <= 1'b0;
      gateways_27_waitCompletion <= 1'b0;
      gateways_28_ip <= 1'b0;
      gateways_28_waitCompletion <= 1'b0;
      gateways_29_ip <= 1'b0;
      gateways_29_waitCompletion <= 1'b0;
      gateways_30_ip <= 1'b0;
      gateways_30_waitCompletion <= 1'b0;
      gateways_0_priority_driver <= 2'b00;
      gateways_1_priority_driver <= 2'b00;
      gateways_2_priority_driver <= 2'b00;
      gateways_3_priority_driver <= 2'b00;
      gateways_4_priority_driver <= 2'b00;
      gateways_5_priority_driver <= 2'b00;
      gateways_6_priority_driver <= 2'b00;
      gateways_7_priority_driver <= 2'b00;
      gateways_8_priority_driver <= 2'b00;
      gateways_9_priority_driver <= 2'b00;
      gateways_10_priority_driver <= 2'b00;
      gateways_11_priority_driver <= 2'b00;
      gateways_12_priority_driver <= 2'b00;
      gateways_13_priority_driver <= 2'b00;
      gateways_14_priority_driver <= 2'b00;
      gateways_15_priority_driver <= 2'b00;
      gateways_16_priority_driver <= 2'b00;
      gateways_17_priority_driver <= 2'b00;
      gateways_18_priority_driver <= 2'b00;
      gateways_19_priority_driver <= 2'b00;
      gateways_20_priority_driver <= 2'b00;
      gateways_21_priority_driver <= 2'b00;
      gateways_22_priority_driver <= 2'b00;
      gateways_23_priority_driver <= 2'b00;
      gateways_24_priority_driver <= 2'b00;
      gateways_25_priority_driver <= 2'b00;
      gateways_26_priority_driver <= 2'b00;
      gateways_27_priority_driver <= 2'b00;
      gateways_28_priority_driver <= 2'b00;
      gateways_29_priority_driver <= 2'b00;
      gateways_30_priority_driver <= 2'b00;
      mapping_coherencyStall_value <= 1'b0;
      targets_0_threshold_driver <= 2'b00;
      targets_0_ie_0_driver <= 1'b0;
      targets_0_ie_1_driver <= 1'b0;
      targets_0_ie_2_driver <= 1'b0;
      targets_0_ie_3_driver <= 1'b0;
      targets_0_ie_4_driver <= 1'b0;
      targets_0_ie_5_driver <= 1'b0;
      targets_0_ie_6_driver <= 1'b0;
      targets_0_ie_7_driver <= 1'b0;
      targets_0_ie_8_driver <= 1'b0;
      targets_0_ie_9_driver <= 1'b0;
      targets_0_ie_10_driver <= 1'b0;
      targets_0_ie_11_driver <= 1'b0;
      targets_0_ie_12_driver <= 1'b0;
      targets_0_ie_13_driver <= 1'b0;
      targets_0_ie_14_driver <= 1'b0;
      targets_0_ie_15_driver <= 1'b0;
      targets_0_ie_16_driver <= 1'b0;
      targets_0_ie_17_driver <= 1'b0;
      targets_0_ie_18_driver <= 1'b0;
      targets_0_ie_19_driver <= 1'b0;
      targets_0_ie_20_driver <= 1'b0;
      targets_0_ie_21_driver <= 1'b0;
      targets_0_ie_22_driver <= 1'b0;
      targets_0_ie_23_driver <= 1'b0;
      targets_0_ie_24_driver <= 1'b0;
      targets_0_ie_25_driver <= 1'b0;
      targets_0_ie_26_driver <= 1'b0;
      targets_0_ie_27_driver <= 1'b0;
      targets_0_ie_28_driver <= 1'b0;
      targets_0_ie_29_driver <= 1'b0;
      targets_0_ie_30_driver <= 1'b0;
      targets_1_threshold_driver <= 2'b00;
      targets_1_ie_0_driver <= 1'b0;
      targets_1_ie_1_driver <= 1'b0;
      targets_1_ie_2_driver <= 1'b0;
      targets_1_ie_3_driver <= 1'b0;
      targets_1_ie_4_driver <= 1'b0;
      targets_1_ie_5_driver <= 1'b0;
      targets_1_ie_6_driver <= 1'b0;
      targets_1_ie_7_driver <= 1'b0;
      targets_1_ie_8_driver <= 1'b0;
      targets_1_ie_9_driver <= 1'b0;
      targets_1_ie_10_driver <= 1'b0;
      targets_1_ie_11_driver <= 1'b0;
      targets_1_ie_12_driver <= 1'b0;
      targets_1_ie_13_driver <= 1'b0;
      targets_1_ie_14_driver <= 1'b0;
      targets_1_ie_15_driver <= 1'b0;
      targets_1_ie_16_driver <= 1'b0;
      targets_1_ie_17_driver <= 1'b0;
      targets_1_ie_18_driver <= 1'b0;
      targets_1_ie_19_driver <= 1'b0;
      targets_1_ie_20_driver <= 1'b0;
      targets_1_ie_21_driver <= 1'b0;
      targets_1_ie_22_driver <= 1'b0;
      targets_1_ie_23_driver <= 1'b0;
      targets_1_ie_24_driver <= 1'b0;
      targets_1_ie_25_driver <= 1'b0;
      targets_1_ie_26_driver <= 1'b0;
      targets_1_ie_27_driver <= 1'b0;
      targets_1_ie_28_driver <= 1'b0;
      targets_1_ie_29_driver <= 1'b0;
      targets_1_ie_30_driver <= 1'b0;
      factory_rspAsync_rValid <= 1'b0;
    end else begin
      if(when_PlicGateway_l21) begin
        gateways_0_ip <= _zz_gateways_0_ip;
        gateways_0_waitCompletion <= _zz_gateways_0_ip;
      end
      if(when_PlicGateway_l21_1) begin
        gateways_1_ip <= _zz_gateways_1_ip;
        gateways_1_waitCompletion <= _zz_gateways_1_ip;
      end
      if(when_PlicGateway_l21_2) begin
        gateways_2_ip <= _zz_gateways_2_ip;
        gateways_2_waitCompletion <= _zz_gateways_2_ip;
      end
      if(when_PlicGateway_l21_3) begin
        gateways_3_ip <= _zz_gateways_3_ip;
        gateways_3_waitCompletion <= _zz_gateways_3_ip;
      end
      if(when_PlicGateway_l21_4) begin
        gateways_4_ip <= _zz_gateways_4_ip;
        gateways_4_waitCompletion <= _zz_gateways_4_ip;
      end
      if(when_PlicGateway_l21_5) begin
        gateways_5_ip <= _zz_gateways_5_ip;
        gateways_5_waitCompletion <= _zz_gateways_5_ip;
      end
      if(when_PlicGateway_l21_6) begin
        gateways_6_ip <= _zz_gateways_6_ip;
        gateways_6_waitCompletion <= _zz_gateways_6_ip;
      end
      if(when_PlicGateway_l21_7) begin
        gateways_7_ip <= _zz_gateways_7_ip;
        gateways_7_waitCompletion <= _zz_gateways_7_ip;
      end
      if(when_PlicGateway_l21_8) begin
        gateways_8_ip <= _zz_gateways_8_ip;
        gateways_8_waitCompletion <= _zz_gateways_8_ip;
      end
      if(when_PlicGateway_l21_9) begin
        gateways_9_ip <= _zz_gateways_9_ip;
        gateways_9_waitCompletion <= _zz_gateways_9_ip;
      end
      if(when_PlicGateway_l21_10) begin
        gateways_10_ip <= _zz_gateways_10_ip;
        gateways_10_waitCompletion <= _zz_gateways_10_ip;
      end
      if(when_PlicGateway_l21_11) begin
        gateways_11_ip <= _zz_gateways_11_ip;
        gateways_11_waitCompletion <= _zz_gateways_11_ip;
      end
      if(when_PlicGateway_l21_12) begin
        gateways_12_ip <= _zz_gateways_12_ip;
        gateways_12_waitCompletion <= _zz_gateways_12_ip;
      end
      if(when_PlicGateway_l21_13) begin
        gateways_13_ip <= _zz_gateways_13_ip;
        gateways_13_waitCompletion <= _zz_gateways_13_ip;
      end
      if(when_PlicGateway_l21_14) begin
        gateways_14_ip <= _zz_gateways_14_ip;
        gateways_14_waitCompletion <= _zz_gateways_14_ip;
      end
      if(when_PlicGateway_l21_15) begin
        gateways_15_ip <= _zz_gateways_15_ip;
        gateways_15_waitCompletion <= _zz_gateways_15_ip;
      end
      if(when_PlicGateway_l21_16) begin
        gateways_16_ip <= _zz_gateways_16_ip;
        gateways_16_waitCompletion <= _zz_gateways_16_ip;
      end
      if(when_PlicGateway_l21_17) begin
        gateways_17_ip <= _zz_gateways_17_ip;
        gateways_17_waitCompletion <= _zz_gateways_17_ip;
      end
      if(when_PlicGateway_l21_18) begin
        gateways_18_ip <= _zz_gateways_18_ip;
        gateways_18_waitCompletion <= _zz_gateways_18_ip;
      end
      if(when_PlicGateway_l21_19) begin
        gateways_19_ip <= _zz_gateways_19_ip;
        gateways_19_waitCompletion <= _zz_gateways_19_ip;
      end
      if(when_PlicGateway_l21_20) begin
        gateways_20_ip <= _zz_gateways_20_ip;
        gateways_20_waitCompletion <= _zz_gateways_20_ip;
      end
      if(when_PlicGateway_l21_21) begin
        gateways_21_ip <= _zz_gateways_21_ip;
        gateways_21_waitCompletion <= _zz_gateways_21_ip;
      end
      if(when_PlicGateway_l21_22) begin
        gateways_22_ip <= _zz_gateways_22_ip;
        gateways_22_waitCompletion <= _zz_gateways_22_ip;
      end
      if(when_PlicGateway_l21_23) begin
        gateways_23_ip <= _zz_gateways_23_ip;
        gateways_23_waitCompletion <= _zz_gateways_23_ip;
      end
      if(when_PlicGateway_l21_24) begin
        gateways_24_ip <= _zz_gateways_24_ip;
        gateways_24_waitCompletion <= _zz_gateways_24_ip;
      end
      if(when_PlicGateway_l21_25) begin
        gateways_25_ip <= _zz_gateways_25_ip;
        gateways_25_waitCompletion <= _zz_gateways_25_ip;
      end
      if(when_PlicGateway_l21_26) begin
        gateways_26_ip <= _zz_gateways_26_ip;
        gateways_26_waitCompletion <= _zz_gateways_26_ip;
      end
      if(when_PlicGateway_l21_27) begin
        gateways_27_ip <= _zz_gateways_27_ip;
        gateways_27_waitCompletion <= _zz_gateways_27_ip;
      end
      if(when_PlicGateway_l21_28) begin
        gateways_28_ip <= _zz_gateways_28_ip;
        gateways_28_waitCompletion <= _zz_gateways_28_ip;
      end
      if(when_PlicGateway_l21_29) begin
        gateways_29_ip <= _zz_gateways_29_ip;
        gateways_29_waitCompletion <= _zz_gateways_29_ip;
      end
      if(when_PlicGateway_l21_30) begin
        gateways_30_ip <= _zz_gateways_30_ip;
        gateways_30_waitCompletion <= _zz_gateways_30_ip;
      end
      if(mapping_claim_valid) begin
        case(mapping_claim_payload)
          5'h01 : begin
            gateways_0_ip <= 1'b0;
          end
          5'h02 : begin
            gateways_1_ip <= 1'b0;
          end
          5'h03 : begin
            gateways_2_ip <= 1'b0;
          end
          5'h04 : begin
            gateways_3_ip <= 1'b0;
          end
          5'h05 : begin
            gateways_4_ip <= 1'b0;
          end
          5'h06 : begin
            gateways_5_ip <= 1'b0;
          end
          5'h07 : begin
            gateways_6_ip <= 1'b0;
          end
          5'h08 : begin
            gateways_7_ip <= 1'b0;
          end
          5'h09 : begin
            gateways_8_ip <= 1'b0;
          end
          5'h0a : begin
            gateways_9_ip <= 1'b0;
          end
          5'h0b : begin
            gateways_10_ip <= 1'b0;
          end
          5'h0c : begin
            gateways_11_ip <= 1'b0;
          end
          5'h0d : begin
            gateways_12_ip <= 1'b0;
          end
          5'h0e : begin
            gateways_13_ip <= 1'b0;
          end
          5'h0f : begin
            gateways_14_ip <= 1'b0;
          end
          5'h10 : begin
            gateways_15_ip <= 1'b0;
          end
          5'h11 : begin
            gateways_16_ip <= 1'b0;
          end
          5'h12 : begin
            gateways_17_ip <= 1'b0;
          end
          5'h13 : begin
            gateways_18_ip <= 1'b0;
          end
          5'h14 : begin
            gateways_19_ip <= 1'b0;
          end
          5'h15 : begin
            gateways_20_ip <= 1'b0;
          end
          5'h16 : begin
            gateways_21_ip <= 1'b0;
          end
          5'h17 : begin
            gateways_22_ip <= 1'b0;
          end
          5'h18 : begin
            gateways_23_ip <= 1'b0;
          end
          5'h19 : begin
            gateways_24_ip <= 1'b0;
          end
          5'h1a : begin
            gateways_25_ip <= 1'b0;
          end
          5'h1b : begin
            gateways_26_ip <= 1'b0;
          end
          5'h1c : begin
            gateways_27_ip <= 1'b0;
          end
          5'h1d : begin
            gateways_28_ip <= 1'b0;
          end
          5'h1e : begin
            gateways_29_ip <= 1'b0;
          end
          5'h1f : begin
            gateways_30_ip <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      if(mapping_completion_valid) begin
        case(mapping_completion_payload)
          5'h01 : begin
            gateways_0_waitCompletion <= 1'b0;
          end
          5'h02 : begin
            gateways_1_waitCompletion <= 1'b0;
          end
          5'h03 : begin
            gateways_2_waitCompletion <= 1'b0;
          end
          5'h04 : begin
            gateways_3_waitCompletion <= 1'b0;
          end
          5'h05 : begin
            gateways_4_waitCompletion <= 1'b0;
          end
          5'h06 : begin
            gateways_5_waitCompletion <= 1'b0;
          end
          5'h07 : begin
            gateways_6_waitCompletion <= 1'b0;
          end
          5'h08 : begin
            gateways_7_waitCompletion <= 1'b0;
          end
          5'h09 : begin
            gateways_8_waitCompletion <= 1'b0;
          end
          5'h0a : begin
            gateways_9_waitCompletion <= 1'b0;
          end
          5'h0b : begin
            gateways_10_waitCompletion <= 1'b0;
          end
          5'h0c : begin
            gateways_11_waitCompletion <= 1'b0;
          end
          5'h0d : begin
            gateways_12_waitCompletion <= 1'b0;
          end
          5'h0e : begin
            gateways_13_waitCompletion <= 1'b0;
          end
          5'h0f : begin
            gateways_14_waitCompletion <= 1'b0;
          end
          5'h10 : begin
            gateways_15_waitCompletion <= 1'b0;
          end
          5'h11 : begin
            gateways_16_waitCompletion <= 1'b0;
          end
          5'h12 : begin
            gateways_17_waitCompletion <= 1'b0;
          end
          5'h13 : begin
            gateways_18_waitCompletion <= 1'b0;
          end
          5'h14 : begin
            gateways_19_waitCompletion <= 1'b0;
          end
          5'h15 : begin
            gateways_20_waitCompletion <= 1'b0;
          end
          5'h16 : begin
            gateways_21_waitCompletion <= 1'b0;
          end
          5'h17 : begin
            gateways_22_waitCompletion <= 1'b0;
          end
          5'h18 : begin
            gateways_23_waitCompletion <= 1'b0;
          end
          5'h19 : begin
            gateways_24_waitCompletion <= 1'b0;
          end
          5'h1a : begin
            gateways_25_waitCompletion <= 1'b0;
          end
          5'h1b : begin
            gateways_26_waitCompletion <= 1'b0;
          end
          5'h1c : begin
            gateways_27_waitCompletion <= 1'b0;
          end
          5'h1d : begin
            gateways_28_waitCompletion <= 1'b0;
          end
          5'h1e : begin
            gateways_29_waitCompletion <= 1'b0;
          end
          5'h1f : begin
            gateways_30_waitCompletion <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      mapping_coherencyStall_value <= mapping_coherencyStall_valueNext;
      if(factory_rspAsync_ready) begin
        factory_rspAsync_rValid <= factory_rspAsync_valid;
      end
      case(factory_address)
        22'h000004 : begin
          if(factory_doWrite) begin
            gateways_0_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000008 : begin
          if(factory_doWrite) begin
            gateways_1_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h00000c : begin
          if(factory_doWrite) begin
            gateways_2_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000010 : begin
          if(factory_doWrite) begin
            gateways_3_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000014 : begin
          if(factory_doWrite) begin
            gateways_4_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000018 : begin
          if(factory_doWrite) begin
            gateways_5_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h00001c : begin
          if(factory_doWrite) begin
            gateways_6_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000020 : begin
          if(factory_doWrite) begin
            gateways_7_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000024 : begin
          if(factory_doWrite) begin
            gateways_8_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000028 : begin
          if(factory_doWrite) begin
            gateways_9_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h00002c : begin
          if(factory_doWrite) begin
            gateways_10_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000030 : begin
          if(factory_doWrite) begin
            gateways_11_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000034 : begin
          if(factory_doWrite) begin
            gateways_12_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000038 : begin
          if(factory_doWrite) begin
            gateways_13_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h00003c : begin
          if(factory_doWrite) begin
            gateways_14_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000040 : begin
          if(factory_doWrite) begin
            gateways_15_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000044 : begin
          if(factory_doWrite) begin
            gateways_16_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000048 : begin
          if(factory_doWrite) begin
            gateways_17_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h00004c : begin
          if(factory_doWrite) begin
            gateways_18_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000050 : begin
          if(factory_doWrite) begin
            gateways_19_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000054 : begin
          if(factory_doWrite) begin
            gateways_20_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000058 : begin
          if(factory_doWrite) begin
            gateways_21_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h00005c : begin
          if(factory_doWrite) begin
            gateways_22_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000060 : begin
          if(factory_doWrite) begin
            gateways_23_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000064 : begin
          if(factory_doWrite) begin
            gateways_24_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000068 : begin
          if(factory_doWrite) begin
            gateways_25_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h00006c : begin
          if(factory_doWrite) begin
            gateways_26_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000070 : begin
          if(factory_doWrite) begin
            gateways_27_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000074 : begin
          if(factory_doWrite) begin
            gateways_28_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h000078 : begin
          if(factory_doWrite) begin
            gateways_29_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h00007c : begin
          if(factory_doWrite) begin
            gateways_30_priority_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h200000 : begin
          if(factory_doWrite) begin
            targets_0_threshold_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h002000 : begin
          if(factory_doWrite) begin
            targets_0_ie_0_driver <= io_bus_a_payload_data[1];
            targets_0_ie_1_driver <= io_bus_a_payload_data[2];
            targets_0_ie_2_driver <= io_bus_a_payload_data[3];
            targets_0_ie_3_driver <= io_bus_a_payload_data[4];
            targets_0_ie_4_driver <= io_bus_a_payload_data[5];
            targets_0_ie_5_driver <= io_bus_a_payload_data[6];
            targets_0_ie_6_driver <= io_bus_a_payload_data[7];
            targets_0_ie_7_driver <= io_bus_a_payload_data[8];
            targets_0_ie_8_driver <= io_bus_a_payload_data[9];
            targets_0_ie_9_driver <= io_bus_a_payload_data[10];
            targets_0_ie_10_driver <= io_bus_a_payload_data[11];
            targets_0_ie_11_driver <= io_bus_a_payload_data[12];
            targets_0_ie_12_driver <= io_bus_a_payload_data[13];
            targets_0_ie_13_driver <= io_bus_a_payload_data[14];
            targets_0_ie_14_driver <= io_bus_a_payload_data[15];
            targets_0_ie_15_driver <= io_bus_a_payload_data[16];
            targets_0_ie_16_driver <= io_bus_a_payload_data[17];
            targets_0_ie_17_driver <= io_bus_a_payload_data[18];
            targets_0_ie_18_driver <= io_bus_a_payload_data[19];
            targets_0_ie_19_driver <= io_bus_a_payload_data[20];
            targets_0_ie_20_driver <= io_bus_a_payload_data[21];
            targets_0_ie_21_driver <= io_bus_a_payload_data[22];
            targets_0_ie_22_driver <= io_bus_a_payload_data[23];
            targets_0_ie_23_driver <= io_bus_a_payload_data[24];
            targets_0_ie_24_driver <= io_bus_a_payload_data[25];
            targets_0_ie_25_driver <= io_bus_a_payload_data[26];
            targets_0_ie_26_driver <= io_bus_a_payload_data[27];
            targets_0_ie_27_driver <= io_bus_a_payload_data[28];
            targets_0_ie_28_driver <= io_bus_a_payload_data[29];
            targets_0_ie_29_driver <= io_bus_a_payload_data[30];
            targets_0_ie_30_driver <= io_bus_a_payload_data[31];
          end
        end
        22'h201000 : begin
          if(factory_doWrite) begin
            targets_1_threshold_driver <= io_bus_a_payload_data[1 : 0];
          end
        end
        22'h002080 : begin
          if(factory_doWrite) begin
            targets_1_ie_0_driver <= io_bus_a_payload_data[1];
            targets_1_ie_1_driver <= io_bus_a_payload_data[2];
            targets_1_ie_2_driver <= io_bus_a_payload_data[3];
            targets_1_ie_3_driver <= io_bus_a_payload_data[4];
            targets_1_ie_4_driver <= io_bus_a_payload_data[5];
            targets_1_ie_5_driver <= io_bus_a_payload_data[6];
            targets_1_ie_6_driver <= io_bus_a_payload_data[7];
            targets_1_ie_7_driver <= io_bus_a_payload_data[8];
            targets_1_ie_8_driver <= io_bus_a_payload_data[9];
            targets_1_ie_9_driver <= io_bus_a_payload_data[10];
            targets_1_ie_10_driver <= io_bus_a_payload_data[11];
            targets_1_ie_11_driver <= io_bus_a_payload_data[12];
            targets_1_ie_12_driver <= io_bus_a_payload_data[13];
            targets_1_ie_13_driver <= io_bus_a_payload_data[14];
            targets_1_ie_14_driver <= io_bus_a_payload_data[15];
            targets_1_ie_15_driver <= io_bus_a_payload_data[16];
            targets_1_ie_16_driver <= io_bus_a_payload_data[17];
            targets_1_ie_17_driver <= io_bus_a_payload_data[18];
            targets_1_ie_18_driver <= io_bus_a_payload_data[19];
            targets_1_ie_19_driver <= io_bus_a_payload_data[20];
            targets_1_ie_20_driver <= io_bus_a_payload_data[21];
            targets_1_ie_21_driver <= io_bus_a_payload_data[22];
            targets_1_ie_22_driver <= io_bus_a_payload_data[23];
            targets_1_ie_23_driver <= io_bus_a_payload_data[24];
            targets_1_ie_24_driver <= io_bus_a_payload_data[25];
            targets_1_ie_25_driver <= io_bus_a_payload_data[26];
            targets_1_ie_26_driver <= io_bus_a_payload_data[27];
            targets_1_ie_27_driver <= io_bus_a_payload_data[28];
            targets_1_ie_28_driver <= io_bus_a_payload_data[29];
            targets_1_ie_29_driver <= io_bus_a_payload_data[30];
            targets_1_ie_30_driver <= io_bus_a_payload_data[31];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge litex_clk) begin
    targets_0_bestRequest_priority <= (_zz_targets_0_bestRequest_priority_6 ? _zz_targets_0_bestRequest_priority_4 : _zz_targets_0_bestRequest_priority_5);
    targets_0_bestRequest_id <= (_zz_targets_0_bestRequest_priority_6 ? (_zz_targets_0_bestRequest_id_80 ? (_zz_targets_0_bestRequest_id_72 ? (_zz_targets_0_bestRequest_id_48 ? _zz_targets_0_bestRequest_id_82 : _zz_targets_0_bestRequest_id_83) : (_zz_targets_0_bestRequest_id_51 ? _zz_targets_0_bestRequest_id_84 : _zz_targets_0_bestRequest_id_85)) : (_zz_targets_0_bestRequest_id_74 ? (_zz_targets_0_bestRequest_id_54 ? _zz_targets_0_bestRequest_id_86 : _zz_targets_0_bestRequest_id_87) : (_zz_targets_0_bestRequest_id_57 ? _zz_targets_0_bestRequest_id_88 : _zz_targets_0_bestRequest_id_89))) : (_zz_targets_0_bestRequest_id_81 ? (_zz_targets_0_bestRequest_id_76 ? (_zz_targets_0_bestRequest_id_60 ? _zz_targets_0_bestRequest_id_90 : _zz_targets_0_bestRequest_id_91) : (_zz_targets_0_bestRequest_id_63 ? _zz_targets_0_bestRequest_id_92 : _zz_targets_0_bestRequest_id_93)) : (_zz_targets_0_bestRequest_id_78 ? (_zz_targets_0_bestRequest_id_66 ? _zz_targets_0_bestRequest_id_94 : _zz_targets_0_bestRequest_id_95) : (_zz_targets_0_bestRequest_id_69 ? _zz_targets_0_bestRequest_id_96 : _zz_targets_0_bestRequest_id_97))));
    targets_0_bestRequest_valid <= (_zz_targets_0_bestRequest_priority_6 ? _zz_targets_0_bestRequest_valid : _zz_targets_0_bestRequest_valid_1);
    targets_1_bestRequest_priority <= (_zz_targets_1_bestRequest_priority_6 ? _zz_targets_1_bestRequest_priority_4 : _zz_targets_1_bestRequest_priority_5);
    targets_1_bestRequest_id <= (_zz_targets_1_bestRequest_priority_6 ? (_zz_targets_1_bestRequest_id_80 ? (_zz_targets_1_bestRequest_id_72 ? (_zz_targets_1_bestRequest_id_48 ? _zz_targets_1_bestRequest_id_82 : _zz_targets_1_bestRequest_id_83) : (_zz_targets_1_bestRequest_id_51 ? _zz_targets_1_bestRequest_id_84 : _zz_targets_1_bestRequest_id_85)) : (_zz_targets_1_bestRequest_id_74 ? (_zz_targets_1_bestRequest_id_54 ? _zz_targets_1_bestRequest_id_86 : _zz_targets_1_bestRequest_id_87) : (_zz_targets_1_bestRequest_id_57 ? _zz_targets_1_bestRequest_id_88 : _zz_targets_1_bestRequest_id_89))) : (_zz_targets_1_bestRequest_id_81 ? (_zz_targets_1_bestRequest_id_76 ? (_zz_targets_1_bestRequest_id_60 ? _zz_targets_1_bestRequest_id_90 : _zz_targets_1_bestRequest_id_91) : (_zz_targets_1_bestRequest_id_63 ? _zz_targets_1_bestRequest_id_92 : _zz_targets_1_bestRequest_id_93)) : (_zz_targets_1_bestRequest_id_78 ? (_zz_targets_1_bestRequest_id_66 ? _zz_targets_1_bestRequest_id_94 : _zz_targets_1_bestRequest_id_95) : (_zz_targets_1_bestRequest_id_69 ? _zz_targets_1_bestRequest_id_96 : _zz_targets_1_bestRequest_id_97))));
    targets_1_bestRequest_valid <= (_zz_targets_1_bestRequest_priority_6 ? _zz_targets_1_bestRequest_valid : _zz_targets_1_bestRequest_valid_1);
    if(factory_rspAsync_ready) begin
      factory_rspAsync_rData_opcode <= factory_rspAsync_payload_opcode;
      factory_rspAsync_rData_param <= factory_rspAsync_payload_param;
      factory_rspAsync_rData_source <= factory_rspAsync_payload_source;
      factory_rspAsync_rData_size <= factory_rspAsync_payload_size;
      factory_rspAsync_rData_denied <= factory_rspAsync_payload_denied;
      factory_rspAsync_rData_data <= factory_rspAsync_payload_data;
      factory_rspAsync_rData_corrupt <= factory_rspAsync_payload_corrupt;
    end
  end


endmodule

module TilelinkClint (
  input  wire          io_bus_a_valid,
  output wire          io_bus_a_ready,
  input  wire [2:0]    io_bus_a_payload_opcode,
  input  wire [2:0]    io_bus_a_payload_param,
  input  wire [2:0]    io_bus_a_payload_source,
  input  wire [15:0]   io_bus_a_payload_address,
  input  wire [2:0]    io_bus_a_payload_size,
  input  wire [3:0]    io_bus_a_payload_mask,
  input  wire [31:0]   io_bus_a_payload_data,
  input  wire          io_bus_a_payload_corrupt,
  output wire          io_bus_d_valid,
  input  wire          io_bus_d_ready,
  output wire [2:0]    io_bus_d_payload_opcode,
  output wire [2:0]    io_bus_d_payload_param,
  output wire [2:0]    io_bus_d_payload_source,
  output wire [2:0]    io_bus_d_payload_size,
  output wire          io_bus_d_payload_denied,
  output wire [31:0]   io_bus_d_payload_data,
  output wire          io_bus_d_payload_corrupt,
  output wire [0:0]    io_timerInterrupt,
  output wire [0:0]    io_softwareInterrupt,
  output wire [63:0]   io_time,
  input  wire          io_stop,
  input  wire          litex_clk,
  input  wire          litex_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  reg        [3:0]    _zz_factory_unburstify_last;
  wire       [15:0]   _zz_factory_unburstify_busA_payload_address;
  wire       [5:0]    _zz_factory_unburstify_busA_payload_address_1;
  wire       [13:0]   _zz_factory_address;
  wire                factory_readErrorFlag;
  wire                factory_writeErrorFlag;
  wire                factory_unburstify_isGet;
  reg        [3:0]    factory_unburstify_counter;
  wire                factory_unburstify_last;
  wire                factory_unburstify_busA_valid;
  wire                factory_unburstify_busA_ready;
  wire       [2:0]    factory_unburstify_busA_payload_opcode;
  wire       [2:0]    factory_unburstify_busA_payload_param;
  wire       [2:0]    factory_unburstify_busA_payload_source;
  wire       [15:0]   factory_unburstify_busA_payload_address;
  wire       [2:0]    factory_unburstify_busA_payload_size;
  wire       [3:0]    factory_unburstify_busA_payload_mask;
  wire       [31:0]   factory_unburstify_busA_payload_data;
  wire                factory_unburstify_busA_payload_corrupt;
  wire                factory_unburstify_busA_fire;
  wire                io_bus_a_fire;
  wire                when_SlaveFactory_l70;
  wire                factory_unburstify_withRsp;
  wire                factory_rspAsync_valid;
  reg                 factory_rspAsync_ready;
  wire       [2:0]    factory_rspAsync_payload_opcode;
  wire       [2:0]    factory_rspAsync_payload_param;
  wire       [2:0]    factory_rspAsync_payload_source;
  wire       [2:0]    factory_rspAsync_payload_size;
  wire                factory_rspAsync_payload_denied;
  reg        [31:0]   factory_rspAsync_payload_data;
  wire                factory_rspAsync_payload_corrupt;
  wire                factory_askWrite;
  wire                factory_askRead;
  wire                factory_doWrite;
  wire                factory_doRead;
  wire       [15:0]   factory_address;
  wire                factory_halt;
  reg                 logic_stop;
  reg        [63:0]   logic_time;
  wire                when_Clint_l39;
  reg        [63:0]   logic_harts_0_cmp;
  reg                 logic_harts_0_timerInterrupt;
  reg                 logic_harts_0_softwareInterrupt;
  reg                 when_Clint_l59;
  reg        [31:0]   _zz_factory_rspAsync_payload_data;
  wire       [2:0]    _zz_factory_rspAsync_payload_opcode;
  wire                factory_rspAsync_stage_valid;
  wire                factory_rspAsync_stage_ready;
  wire       [2:0]    factory_rspAsync_stage_payload_opcode;
  wire       [2:0]    factory_rspAsync_stage_payload_param;
  wire       [2:0]    factory_rspAsync_stage_payload_source;
  wire       [2:0]    factory_rspAsync_stage_payload_size;
  wire                factory_rspAsync_stage_payload_denied;
  wire       [31:0]   factory_rspAsync_stage_payload_data;
  wire                factory_rspAsync_stage_payload_corrupt;
  reg                 factory_rspAsync_rValid;
  reg        [2:0]    factory_rspAsync_rData_opcode;
  reg        [2:0]    factory_rspAsync_rData_param;
  reg        [2:0]    factory_rspAsync_rData_source;
  reg        [2:0]    factory_rspAsync_rData_size;
  reg                 factory_rspAsync_rData_denied;
  reg        [31:0]   factory_rspAsync_rData_data;
  reg                 factory_rspAsync_rData_corrupt;
  wire                when_Stream_l399;
  wire                when_SlaveFactory_l134;
  wire                when_SlaveFactory_l134_1;
  `ifndef SYNTHESIS
  reg [127:0] io_bus_a_payload_opcode_string;
  reg [119:0] io_bus_d_payload_opcode_string;
  reg [127:0] factory_unburstify_busA_payload_opcode_string;
  reg [119:0] factory_rspAsync_payload_opcode_string;
  reg [119:0] _zz_factory_rspAsync_payload_opcode_string;
  reg [119:0] factory_rspAsync_stage_payload_opcode_string;
  reg [119:0] factory_rspAsync_rData_opcode_string;
  `endif


  assign _zz_factory_unburstify_busA_payload_address_1 = ({2'd0,factory_unburstify_counter} <<< 2'd2);
  assign _zz_factory_unburstify_busA_payload_address = {10'd0, _zz_factory_unburstify_busA_payload_address_1};
  assign _zz_factory_address = (factory_unburstify_busA_payload_address >>> 2'd2);
  always @(*) begin
    case(io_bus_a_payload_size)
      3'b000 : _zz_factory_unburstify_last = 4'b0000;
      3'b001 : _zz_factory_unburstify_last = 4'b0000;
      3'b010 : _zz_factory_unburstify_last = 4'b0000;
      3'b011 : _zz_factory_unburstify_last = 4'b0001;
      3'b100 : _zz_factory_unburstify_last = 4'b0011;
      3'b101 : _zz_factory_unburstify_last = 4'b0111;
      default : _zz_factory_unburstify_last = 4'b1111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_bus_a_payload_opcode)
      A_PUT_FULL_DATA : io_bus_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_bus_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_bus_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_bus_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_bus_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_bus_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_bus_d_payload_opcode)
      D_ACCESS_ACK : io_bus_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_bus_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_bus_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_bus_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_bus_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_bus_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(factory_unburstify_busA_payload_opcode)
      A_PUT_FULL_DATA : factory_unburstify_busA_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : factory_unburstify_busA_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : factory_unburstify_busA_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : factory_unburstify_busA_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : factory_unburstify_busA_payload_opcode_string = "ACQUIRE_PERM    ";
      default : factory_unburstify_busA_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(factory_rspAsync_payload_opcode)
      D_ACCESS_ACK : factory_rspAsync_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : factory_rspAsync_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : factory_rspAsync_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : factory_rspAsync_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : factory_rspAsync_payload_opcode_string = "RELEASE_ACK    ";
      default : factory_rspAsync_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_factory_rspAsync_payload_opcode)
      D_ACCESS_ACK : _zz_factory_rspAsync_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_factory_rspAsync_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_factory_rspAsync_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_factory_rspAsync_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_factory_rspAsync_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_factory_rspAsync_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(factory_rspAsync_stage_payload_opcode)
      D_ACCESS_ACK : factory_rspAsync_stage_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : factory_rspAsync_stage_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : factory_rspAsync_stage_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : factory_rspAsync_stage_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : factory_rspAsync_stage_payload_opcode_string = "RELEASE_ACK    ";
      default : factory_rspAsync_stage_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(factory_rspAsync_rData_opcode)
      D_ACCESS_ACK : factory_rspAsync_rData_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : factory_rspAsync_rData_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : factory_rspAsync_rData_opcode_string = "GRANT          ";
      D_GRANT_DATA : factory_rspAsync_rData_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : factory_rspAsync_rData_opcode_string = "RELEASE_ACK    ";
      default : factory_rspAsync_rData_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign factory_readErrorFlag = 1'b0;
  assign factory_writeErrorFlag = 1'b0;
  assign factory_unburstify_isGet = (io_bus_a_payload_opcode == A_GET);
  assign factory_unburstify_last = (factory_unburstify_counter == _zz_factory_unburstify_last);
  assign factory_unburstify_busA_valid = io_bus_a_valid;
  assign factory_unburstify_busA_payload_opcode = io_bus_a_payload_opcode;
  assign factory_unburstify_busA_payload_param = io_bus_a_payload_param;
  assign factory_unburstify_busA_payload_source = io_bus_a_payload_source;
  assign factory_unburstify_busA_payload_size = io_bus_a_payload_size;
  assign factory_unburstify_busA_payload_mask = io_bus_a_payload_mask;
  assign factory_unburstify_busA_payload_data = io_bus_a_payload_data;
  assign factory_unburstify_busA_payload_corrupt = io_bus_a_payload_corrupt;
  assign io_bus_a_ready = (factory_unburstify_busA_ready && ((! factory_unburstify_isGet) || factory_unburstify_last));
  assign factory_unburstify_busA_fire = (factory_unburstify_busA_valid && factory_unburstify_busA_ready);
  assign io_bus_a_fire = (io_bus_a_valid && io_bus_a_ready);
  assign when_SlaveFactory_l70 = (io_bus_a_fire && (factory_unburstify_isGet || factory_unburstify_last));
  assign factory_unburstify_busA_payload_address = (io_bus_a_payload_address | _zz_factory_unburstify_busA_payload_address);
  assign factory_unburstify_withRsp = (factory_unburstify_isGet || factory_unburstify_last);
  assign factory_askWrite = (factory_unburstify_busA_valid && (|{(factory_unburstify_busA_payload_opcode == A_PUT_PARTIAL_DATA),(factory_unburstify_busA_payload_opcode == A_PUT_FULL_DATA)}));
  assign factory_askRead = (factory_unburstify_busA_valid && (|(factory_unburstify_busA_payload_opcode == A_GET)));
  assign factory_doWrite = (factory_askWrite && factory_unburstify_busA_ready);
  assign factory_doRead = (factory_askRead && factory_unburstify_busA_ready);
  assign factory_address = ({2'd0,_zz_factory_address} <<< 2'd2);
  assign factory_halt = 1'b0;
  always @(*) begin
    logic_stop = 1'b0;
    if(io_stop) begin
      logic_stop = 1'b1;
    end
  end

  assign when_Clint_l39 = (! logic_stop);
  always @(*) begin
    when_Clint_l59 = 1'b0;
    case(factory_address)
      16'hbff8 : begin
        if(factory_doRead) begin
          when_Clint_l59 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign io_timerInterrupt[0] = logic_harts_0_timerInterrupt;
  assign io_softwareInterrupt[0] = logic_harts_0_softwareInterrupt;
  assign io_time = logic_time;
  assign factory_unburstify_busA_ready = (factory_rspAsync_ready && (! factory_halt));
  assign factory_rspAsync_valid = ((factory_unburstify_busA_valid && (! factory_halt)) && factory_unburstify_withRsp);
  always @(*) begin
    factory_rspAsync_payload_data = 32'h0;
    case(factory_address)
      16'hbff8 : begin
        factory_rspAsync_payload_data[31 : 0] = logic_time[31 : 0];
      end
      16'hbffc : begin
        factory_rspAsync_payload_data[31 : 0] = _zz_factory_rspAsync_payload_data;
      end
      16'h0 : begin
        factory_rspAsync_payload_data[0 : 0] = logic_harts_0_softwareInterrupt;
      end
      default : begin
      end
    endcase
  end

  assign _zz_factory_rspAsync_payload_opcode = ((|(factory_unburstify_busA_payload_opcode == A_GET)) ? D_ACCESS_ACK_DATA : D_ACCESS_ACK);
  assign factory_rspAsync_payload_opcode = _zz_factory_rspAsync_payload_opcode;
  assign factory_rspAsync_payload_param = 3'b000;
  assign factory_rspAsync_payload_source = factory_unburstify_busA_payload_source;
  assign factory_rspAsync_payload_size = factory_unburstify_busA_payload_size;
  assign factory_rspAsync_payload_corrupt = 1'b0;
  assign factory_rspAsync_payload_denied = 1'b0;
  always @(*) begin
    factory_rspAsync_ready = factory_rspAsync_stage_ready;
    if(when_Stream_l399) begin
      factory_rspAsync_ready = 1'b1;
    end
  end

  assign when_Stream_l399 = (! factory_rspAsync_stage_valid);
  assign factory_rspAsync_stage_valid = factory_rspAsync_rValid;
  assign factory_rspAsync_stage_payload_opcode = factory_rspAsync_rData_opcode;
  assign factory_rspAsync_stage_payload_param = factory_rspAsync_rData_param;
  assign factory_rspAsync_stage_payload_source = factory_rspAsync_rData_source;
  assign factory_rspAsync_stage_payload_size = factory_rspAsync_rData_size;
  assign factory_rspAsync_stage_payload_denied = factory_rspAsync_rData_denied;
  assign factory_rspAsync_stage_payload_data = factory_rspAsync_rData_data;
  assign factory_rspAsync_stage_payload_corrupt = factory_rspAsync_rData_corrupt;
  assign io_bus_d_valid = factory_rspAsync_stage_valid;
  assign factory_rspAsync_stage_ready = io_bus_d_ready;
  assign io_bus_d_payload_opcode = factory_rspAsync_stage_payload_opcode;
  assign io_bus_d_payload_param = factory_rspAsync_stage_payload_param;
  assign io_bus_d_payload_source = factory_rspAsync_stage_payload_source;
  assign io_bus_d_payload_size = factory_rspAsync_stage_payload_size;
  assign io_bus_d_payload_denied = factory_rspAsync_stage_payload_denied;
  assign io_bus_d_payload_data = factory_rspAsync_stage_payload_data;
  assign io_bus_d_payload_corrupt = factory_rspAsync_stage_payload_corrupt;
  assign when_SlaveFactory_l134 = ((factory_address & (~ 16'h0003)) == 16'h4000);
  assign when_SlaveFactory_l134_1 = ((factory_address & (~ 16'h0003)) == 16'h4004);
  always @(posedge litex_clk or posedge litex_reset) begin
    if(litex_reset) begin
      factory_unburstify_counter <= 4'b0000;
      logic_time <= 64'h0;
      logic_harts_0_softwareInterrupt <= 1'b0;
      factory_rspAsync_rValid <= 1'b0;
    end else begin
      if(factory_unburstify_busA_fire) begin
        factory_unburstify_counter <= (factory_unburstify_counter + 4'b0001);
        if(when_SlaveFactory_l70) begin
          factory_unburstify_counter <= 4'b0000;
        end
      end
      if(when_Clint_l39) begin
        logic_time <= (logic_time + 64'h0000000000000001);
      end
      if(factory_rspAsync_ready) begin
        factory_rspAsync_rValid <= factory_rspAsync_valid;
      end
      case(factory_address)
        16'h0 : begin
          if(factory_doWrite) begin
            logic_harts_0_softwareInterrupt <= factory_unburstify_busA_payload_data[0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge litex_clk) begin
    logic_harts_0_timerInterrupt <= (logic_harts_0_cmp <= logic_time);
    if(when_Clint_l59) begin
      _zz_factory_rspAsync_payload_data <= logic_time[63 : 32];
    end
    if(factory_rspAsync_ready) begin
      factory_rspAsync_rData_opcode <= factory_rspAsync_payload_opcode;
      factory_rspAsync_rData_param <= factory_rspAsync_payload_param;
      factory_rspAsync_rData_source <= factory_rspAsync_payload_source;
      factory_rspAsync_rData_size <= factory_rspAsync_payload_size;
      factory_rspAsync_rData_denied <= factory_rspAsync_payload_denied;
      factory_rspAsync_rData_data <= factory_rspAsync_payload_data;
      factory_rspAsync_rData_corrupt <= factory_rspAsync_payload_corrupt;
    end
    if(when_SlaveFactory_l134) begin
      if(factory_doWrite) begin
        logic_harts_0_cmp[31 : 0] <= factory_unburstify_busA_payload_data[31 : 0];
      end
    end
    if(when_SlaveFactory_l134_1) begin
      if(factory_doWrite) begin
        logic_harts_0_cmp[63 : 32] <= factory_unburstify_busA_payload_data[31 : 0];
      end
    end
  end


endmodule

module Decoder (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [1:0]    io_up_a_payload_source,
  input  wire [31:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [7:0]    io_up_a_payload_mask,
  input  wire [63:0]   io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [1:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [63:0]   io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_downs_0_a_valid,
  input  wire          io_downs_0_a_ready,
  output wire [2:0]    io_downs_0_a_payload_opcode,
  output wire [2:0]    io_downs_0_a_payload_param,
  output wire [1:0]    io_downs_0_a_payload_source,
  output wire [31:0]   io_downs_0_a_payload_address,
  output wire [2:0]    io_downs_0_a_payload_size,
  output wire [7:0]    io_downs_0_a_payload_mask,
  output wire [63:0]   io_downs_0_a_payload_data,
  output wire          io_downs_0_a_payload_corrupt,
  input  wire          io_downs_0_d_valid,
  output wire          io_downs_0_d_ready,
  input  wire [2:0]    io_downs_0_d_payload_opcode,
  input  wire [2:0]    io_downs_0_d_payload_param,
  input  wire [1:0]    io_downs_0_d_payload_source,
  input  wire [2:0]    io_downs_0_d_payload_size,
  input  wire          io_downs_0_d_payload_denied,
  input  wire [63:0]   io_downs_0_d_payload_data,
  input  wire          io_downs_0_d_payload_corrupt,
  output wire          io_downs_1_a_valid,
  input  wire          io_downs_1_a_ready,
  output wire [2:0]    io_downs_1_a_payload_opcode,
  output wire [2:0]    io_downs_1_a_payload_param,
  output wire [1:0]    io_downs_1_a_payload_source,
  output wire [31:0]   io_downs_1_a_payload_address,
  output wire [2:0]    io_downs_1_a_payload_size,
  output wire [7:0]    io_downs_1_a_payload_mask,
  output wire [63:0]   io_downs_1_a_payload_data,
  output wire          io_downs_1_a_payload_corrupt,
  input  wire          io_downs_1_d_valid,
  output wire          io_downs_1_d_ready,
  input  wire [2:0]    io_downs_1_d_payload_opcode,
  input  wire [2:0]    io_downs_1_d_payload_param,
  input  wire [1:0]    io_downs_1_d_payload_source,
  input  wire [2:0]    io_downs_1_d_payload_size,
  input  wire          io_downs_1_d_payload_denied,
  input  wire [63:0]   io_downs_1_d_payload_data,
  input  wire          io_downs_1_d_payload_corrupt,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                d_arbiter_io_inputs_0_ready;
  wire                d_arbiter_io_inputs_1_ready;
  wire                d_arbiter_io_output_valid;
  wire       [2:0]    d_arbiter_io_output_payload_opcode;
  wire       [2:0]    d_arbiter_io_output_payload_param;
  wire       [1:0]    d_arbiter_io_output_payload_source;
  wire       [2:0]    d_arbiter_io_output_payload_size;
  wire                d_arbiter_io_output_payload_denied;
  wire       [63:0]   d_arbiter_io_output_payload_data;
  wire                d_arbiter_io_output_payload_corrupt;
  wire       [0:0]    d_arbiter_io_chosen;
  wire       [1:0]    d_arbiter_io_chosenOH;
  wire       [0:0]    _zz_a_logic_0_hit;
  wire       [0:0]    _zz_a_logic_1_hit;
  reg        [1:0]    _zz_1;
  wire       [1:0]    _zz_2;
  wire                downs_0_a_valid;
  wire                downs_0_a_ready;
  wire       [2:0]    downs_0_a_payload_opcode;
  wire       [2:0]    downs_0_a_payload_param;
  wire       [1:0]    downs_0_a_payload_source;
  wire       [31:0]   downs_0_a_payload_address;
  wire       [2:0]    downs_0_a_payload_size;
  wire       [7:0]    downs_0_a_payload_mask;
  wire       [63:0]   downs_0_a_payload_data;
  wire                downs_0_a_payload_corrupt;
  wire                downs_0_d_valid;
  wire                downs_0_d_ready;
  wire       [2:0]    downs_0_d_payload_opcode;
  wire       [2:0]    downs_0_d_payload_param;
  wire       [1:0]    downs_0_d_payload_source;
  wire       [2:0]    downs_0_d_payload_size;
  wire                downs_0_d_payload_denied;
  wire       [63:0]   downs_0_d_payload_data;
  wire                downs_0_d_payload_corrupt;
  wire                downs_1_a_valid;
  wire                downs_1_a_ready;
  wire       [2:0]    downs_1_a_payload_opcode;
  wire       [2:0]    downs_1_a_payload_param;
  wire       [1:0]    downs_1_a_payload_source;
  wire       [31:0]   downs_1_a_payload_address;
  wire       [2:0]    downs_1_a_payload_size;
  wire       [7:0]    downs_1_a_payload_mask;
  wire       [63:0]   downs_1_a_payload_data;
  wire                downs_1_a_payload_corrupt;
  wire                downs_1_d_valid;
  wire                downs_1_d_ready;
  wire       [2:0]    downs_1_d_payload_opcode;
  wire       [2:0]    downs_1_d_payload_param;
  wire       [1:0]    downs_1_d_payload_source;
  wire       [2:0]    downs_1_d_payload_size;
  wire                downs_1_d_payload_denied;
  wire       [63:0]   downs_1_d_payload_data;
  wire                downs_1_d_payload_corrupt;
  wire       [34:0]   a_key;
  wire                a_logic_0_hit;
  wire                a_logic_1_hit;
  wire                a_miss;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] io_downs_0_a_payload_opcode_string;
  reg [119:0] io_downs_0_d_payload_opcode_string;
  reg [127:0] io_downs_1_a_payload_opcode_string;
  reg [119:0] io_downs_1_d_payload_opcode_string;
  reg [127:0] downs_0_a_payload_opcode_string;
  reg [119:0] downs_0_d_payload_opcode_string;
  reg [127:0] downs_1_a_payload_opcode_string;
  reg [119:0] downs_1_d_payload_opcode_string;
  `endif


  assign _zz_a_logic_0_hit = (|((a_key & 35'h0c0000000) == 35'h040000000));
  assign _zz_a_logic_1_hit = (|{((a_key & 35'h080000000) == 35'h080000000),((a_key & 35'h040000000) == 35'h0)});
  assign _zz_2 = {io_downs_1_a_valid,io_downs_0_a_valid};
  StreamArbiter_8 d_arbiter (
    .io_inputs_0_valid           (downs_0_d_valid                        ), //i
    .io_inputs_0_ready           (d_arbiter_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_opcode  (downs_0_d_payload_opcode[2:0]          ), //i
    .io_inputs_0_payload_param   (downs_0_d_payload_param[2:0]           ), //i
    .io_inputs_0_payload_source  (downs_0_d_payload_source[1:0]          ), //i
    .io_inputs_0_payload_size    (downs_0_d_payload_size[2:0]            ), //i
    .io_inputs_0_payload_denied  (downs_0_d_payload_denied               ), //i
    .io_inputs_0_payload_data    (downs_0_d_payload_data[63:0]           ), //i
    .io_inputs_0_payload_corrupt (downs_0_d_payload_corrupt              ), //i
    .io_inputs_1_valid           (downs_1_d_valid                        ), //i
    .io_inputs_1_ready           (d_arbiter_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_opcode  (downs_1_d_payload_opcode[2:0]          ), //i
    .io_inputs_1_payload_param   (downs_1_d_payload_param[2:0]           ), //i
    .io_inputs_1_payload_source  (downs_1_d_payload_source[1:0]          ), //i
    .io_inputs_1_payload_size    (downs_1_d_payload_size[2:0]            ), //i
    .io_inputs_1_payload_denied  (downs_1_d_payload_denied               ), //i
    .io_inputs_1_payload_data    (downs_1_d_payload_data[63:0]           ), //i
    .io_inputs_1_payload_corrupt (downs_1_d_payload_corrupt              ), //i
    .io_output_valid             (d_arbiter_io_output_valid              ), //o
    .io_output_ready             (io_up_d_ready                          ), //i
    .io_output_payload_opcode    (d_arbiter_io_output_payload_opcode[2:0]), //o
    .io_output_payload_param     (d_arbiter_io_output_payload_param[2:0] ), //o
    .io_output_payload_source    (d_arbiter_io_output_payload_source[1:0]), //o
    .io_output_payload_size      (d_arbiter_io_output_payload_size[2:0]  ), //o
    .io_output_payload_denied    (d_arbiter_io_output_payload_denied     ), //o
    .io_output_payload_data      (d_arbiter_io_output_payload_data[63:0] ), //o
    .io_output_payload_corrupt   (d_arbiter_io_output_payload_corrupt    ), //o
    .io_chosen                   (d_arbiter_io_chosen                    ), //o
    .io_chosenOH                 (d_arbiter_io_chosenOH[1:0]             ), //o
    .litex_clk                   (litex_clk                              ), //i
    .cpuResetCtrl_reset          (cpuResetCtrl_reset                     )  //i
  );
  always @(*) begin
    case(_zz_2)
      2'b00 : _zz_1 = 2'b00;
      2'b01 : _zz_1 = 2'b01;
      2'b10 : _zz_1 = 2'b01;
      default : _zz_1 = 2'b10;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_0_a_payload_opcode)
      A_PUT_FULL_DATA : io_downs_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_downs_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_downs_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_downs_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_downs_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_downs_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_0_d_payload_opcode)
      D_ACCESS_ACK : io_downs_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_downs_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_downs_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_downs_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_downs_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_downs_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_1_a_payload_opcode)
      A_PUT_FULL_DATA : io_downs_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_downs_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_downs_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_downs_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_downs_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_downs_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_downs_1_d_payload_opcode)
      D_ACCESS_ACK : io_downs_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_downs_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_downs_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_downs_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_downs_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_downs_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downs_0_a_payload_opcode)
      A_PUT_FULL_DATA : downs_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downs_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downs_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downs_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downs_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : downs_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(downs_0_d_payload_opcode)
      D_ACCESS_ACK : downs_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : downs_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : downs_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : downs_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : downs_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : downs_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(downs_1_a_payload_opcode)
      A_PUT_FULL_DATA : downs_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : downs_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : downs_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : downs_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : downs_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : downs_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(downs_1_d_payload_opcode)
      D_ACCESS_ACK : downs_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : downs_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : downs_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : downs_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : downs_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : downs_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign io_downs_0_a_valid = downs_0_a_valid;
  assign downs_0_a_ready = io_downs_0_a_ready;
  assign io_downs_0_a_payload_opcode = downs_0_a_payload_opcode;
  assign io_downs_0_a_payload_param = downs_0_a_payload_param;
  assign io_downs_0_a_payload_source = downs_0_a_payload_source;
  assign io_downs_0_a_payload_address = downs_0_a_payload_address;
  assign io_downs_0_a_payload_size = downs_0_a_payload_size;
  assign io_downs_0_a_payload_mask = downs_0_a_payload_mask;
  assign io_downs_0_a_payload_data = downs_0_a_payload_data;
  assign io_downs_0_a_payload_corrupt = downs_0_a_payload_corrupt;
  assign downs_0_d_valid = io_downs_0_d_valid;
  assign io_downs_0_d_ready = downs_0_d_ready;
  assign downs_0_d_payload_opcode = io_downs_0_d_payload_opcode;
  assign downs_0_d_payload_param = io_downs_0_d_payload_param;
  assign downs_0_d_payload_source = io_downs_0_d_payload_source;
  assign downs_0_d_payload_size = io_downs_0_d_payload_size;
  assign downs_0_d_payload_denied = io_downs_0_d_payload_denied;
  assign downs_0_d_payload_data = io_downs_0_d_payload_data;
  assign downs_0_d_payload_corrupt = io_downs_0_d_payload_corrupt;
  assign io_downs_1_a_valid = downs_1_a_valid;
  assign downs_1_a_ready = io_downs_1_a_ready;
  assign io_downs_1_a_payload_opcode = downs_1_a_payload_opcode;
  assign io_downs_1_a_payload_param = downs_1_a_payload_param;
  assign io_downs_1_a_payload_source = downs_1_a_payload_source;
  assign io_downs_1_a_payload_address = downs_1_a_payload_address;
  assign io_downs_1_a_payload_size = downs_1_a_payload_size;
  assign io_downs_1_a_payload_mask = downs_1_a_payload_mask;
  assign io_downs_1_a_payload_data = downs_1_a_payload_data;
  assign io_downs_1_a_payload_corrupt = downs_1_a_payload_corrupt;
  assign downs_1_d_valid = io_downs_1_d_valid;
  assign io_downs_1_d_ready = downs_1_d_ready;
  assign downs_1_d_payload_opcode = io_downs_1_d_payload_opcode;
  assign downs_1_d_payload_param = io_downs_1_d_payload_param;
  assign downs_1_d_payload_source = io_downs_1_d_payload_source;
  assign downs_1_d_payload_size = io_downs_1_d_payload_size;
  assign downs_1_d_payload_denied = io_downs_1_d_payload_denied;
  assign downs_1_d_payload_data = io_downs_1_d_payload_data;
  assign downs_1_d_payload_corrupt = io_downs_1_d_payload_corrupt;
  assign a_key = {io_up_a_payload_opcode,io_up_a_payload_address};
  assign a_logic_0_hit = _zz_a_logic_0_hit[0];
  assign downs_0_a_valid = (io_up_a_valid && a_logic_0_hit);
  assign downs_0_a_payload_opcode = io_up_a_payload_opcode;
  assign downs_0_a_payload_param = io_up_a_payload_param;
  assign downs_0_a_payload_source = io_up_a_payload_source;
  assign downs_0_a_payload_mask = io_up_a_payload_mask;
  assign downs_0_a_payload_data = io_up_a_payload_data;
  assign downs_0_a_payload_corrupt = io_up_a_payload_corrupt;
  assign downs_0_a_payload_address = io_up_a_payload_address;
  assign downs_0_a_payload_size = io_up_a_payload_size;
  assign a_logic_1_hit = _zz_a_logic_1_hit[0];
  assign downs_1_a_valid = (io_up_a_valid && a_logic_1_hit);
  assign downs_1_a_payload_opcode = io_up_a_payload_opcode;
  assign downs_1_a_payload_param = io_up_a_payload_param;
  assign downs_1_a_payload_source = io_up_a_payload_source;
  assign downs_1_a_payload_mask = io_up_a_payload_mask;
  assign downs_1_a_payload_data = io_up_a_payload_data;
  assign downs_1_a_payload_corrupt = io_up_a_payload_corrupt;
  assign downs_1_a_payload_address = io_up_a_payload_address;
  assign downs_1_a_payload_size = io_up_a_payload_size;
  assign io_up_a_ready = (|{(downs_1_a_ready && a_logic_1_hit),(downs_0_a_ready && a_logic_0_hit)});
  assign a_miss = (! (|{a_logic_1_hit,a_logic_0_hit}));
  assign downs_0_d_ready = d_arbiter_io_inputs_0_ready;
  assign downs_1_d_ready = d_arbiter_io_inputs_1_ready;
  assign io_up_d_valid = d_arbiter_io_output_valid;
  assign io_up_d_payload_opcode = d_arbiter_io_output_payload_opcode;
  assign io_up_d_payload_param = d_arbiter_io_output_payload_param;
  assign io_up_d_payload_source = d_arbiter_io_output_payload_source;
  assign io_up_d_payload_size = d_arbiter_io_output_payload_size;
  assign io_up_d_payload_denied = d_arbiter_io_output_payload_denied;
  assign io_up_d_payload_data = d_arbiter_io_output_payload_data;
  assign io_up_d_payload_corrupt = d_arbiter_io_output_payload_corrupt;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
    end else begin
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (io_up_a_valid && a_miss))); // Decoder.scala:L106
        `else
          if(!(! (io_up_a_valid && a_miss))) begin
            $display("FAILURE Tilelink decoder miss ???"); // Decoder.scala:L106
            $finish;
          end
        `endif
      `endif
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (io_up_a_valid && (_zz_1 != 2'b01)))); // Decoder.scala:L107
        `else
          if(!(! (io_up_a_valid && (_zz_1 != 2'b01)))) begin
            $display("FAILURE Tilelink decoder miss ???"); // Decoder.scala:L107
            $finish;
          end
        `endif
      `endif
    end
  end


endmodule

module Axi4Bridge (
  input  wire          io_up_a_valid,
  output wire          io_up_a_ready,
  input  wire [2:0]    io_up_a_payload_opcode,
  input  wire [2:0]    io_up_a_payload_param,
  input  wire [1:0]    io_up_a_payload_source,
  input  wire [31:0]   io_up_a_payload_address,
  input  wire [2:0]    io_up_a_payload_size,
  input  wire [15:0]   io_up_a_payload_mask,
  input  wire [127:0]  io_up_a_payload_data,
  input  wire          io_up_a_payload_corrupt,
  output wire          io_up_d_valid,
  input  wire          io_up_d_ready,
  output wire [2:0]    io_up_d_payload_opcode,
  output wire [2:0]    io_up_d_payload_param,
  output wire [1:0]    io_up_d_payload_source,
  output wire [2:0]    io_up_d_payload_size,
  output wire          io_up_d_payload_denied,
  output wire [127:0]  io_up_d_payload_data,
  output wire          io_up_d_payload_corrupt,
  output wire          io_down_aw_valid,
  input  wire          io_down_aw_ready,
  output wire [31:0]   io_down_aw_payload_addr,
  output wire [1:0]    io_down_aw_payload_id,
  output wire [7:0]    io_down_aw_payload_len,
  output wire [2:0]    io_down_aw_payload_size,
  output wire [1:0]    io_down_aw_payload_burst,
  output wire          io_down_aw_payload_allStrb,
  output wire          io_down_w_valid,
  input  wire          io_down_w_ready,
  output wire [127:0]  io_down_w_payload_data,
  output wire [15:0]   io_down_w_payload_strb,
  output wire          io_down_w_payload_last,
  input  wire          io_down_b_valid,
  output wire          io_down_b_ready,
  input  wire [1:0]    io_down_b_payload_id,
  input  wire [1:0]    io_down_b_payload_resp,
  output wire          io_down_ar_valid,
  input  wire          io_down_ar_ready,
  output wire [31:0]   io_down_ar_payload_addr,
  output wire [1:0]    io_down_ar_payload_id,
  output wire [7:0]    io_down_ar_payload_len,
  output wire [2:0]    io_down_ar_payload_size,
  output wire [1:0]    io_down_ar_payload_burst,
  input  wire          io_down_r_valid,
  output wire          io_down_r_ready,
  input  wire [127:0]  io_down_r_payload_data,
  input  wire [1:0]    io_down_r_payload_id,
  input  wire [1:0]    io_down_r_payload_resp,
  input  wire          io_down_r_payload_last,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                a_ctx_io_add_valid;
  wire                a_ctx_io_remove_valid;
  wire                d_arbiter_io_inputs_0_payload_denied;
  wire                d_arbiter_io_inputs_1_payload_denied;
  wire                a_ctx_io_add_ready;
  wire       [2:0]    a_ctx_io_query_context;
  wire                d_arbiter_io_inputs_0_ready;
  wire                d_arbiter_io_inputs_1_ready;
  wire                d_arbiter_io_output_valid;
  wire       [1:0]    d_arbiter_io_output_payload_source;
  wire                d_arbiter_io_output_payload_denied;
  wire                d_arbiter_io_output_payload_last;
  wire       [0:0]    d_arbiter_io_chosen;
  wire       [1:0]    d_arbiter_io_chosenOH;
  reg        [1:0]    _zz_io_up_a_tracker_last;
  reg        [1:0]    _zz_io_up_d_tracker_last;
  reg        [1:0]    _zz_a_cmdFork_tracker_last;
  reg        [1:0]    _zz_a_cmd_len;
  reg        [2:0]    _zz_a_cmd_sizePerBeat;
  reg        [1:0]    _zz_a_data_buffer_tracker_last;
  reg                 a_ctxFull;
  wire                _zz_io_up_a_ready;
  wire                a_halted_valid;
  reg                 a_halted_ready;
  wire       [2:0]    a_halted_payload_opcode;
  wire       [2:0]    a_halted_payload_param;
  wire       [1:0]    a_halted_payload_source;
  wire       [31:0]   a_halted_payload_address;
  wire       [2:0]    a_halted_payload_size;
  wire       [15:0]   a_halted_payload_mask;
  wire       [127:0]  a_halted_payload_data;
  wire                a_halted_payload_corrupt;
  wire                io_up_a_fire;
  reg        [1:0]    io_up_a_tracker_beat;
  wire                io_up_a_tracker_last;
  wire                when_ContextBuffer_l19;
  wire                io_up_d_fire;
  reg        [1:0]    io_up_d_tracker_beat;
  wire                io_up_d_tracker_last;
  wire                a_cmdFork_valid;
  reg                 a_cmdFork_ready;
  wire       [2:0]    a_cmdFork_payload_opcode;
  wire       [2:0]    a_cmdFork_payload_param;
  wire       [1:0]    a_cmdFork_payload_source;
  wire       [31:0]   a_cmdFork_payload_address;
  wire       [2:0]    a_cmdFork_payload_size;
  wire       [15:0]   a_cmdFork_payload_mask;
  wire       [127:0]  a_cmdFork_payload_data;
  wire                a_cmdFork_payload_corrupt;
  wire                a_dataFork_valid;
  reg                 a_dataFork_ready;
  wire       [2:0]    a_dataFork_payload_opcode;
  wire       [2:0]    a_dataFork_payload_param;
  wire       [1:0]    a_dataFork_payload_source;
  wire       [31:0]   a_dataFork_payload_address;
  wire       [2:0]    a_dataFork_payload_size;
  wire       [15:0]   a_dataFork_payload_mask;
  wire       [127:0]  a_dataFork_payload_data;
  wire                a_dataFork_payload_corrupt;
  reg                 a_halted_fork2_logic_linkEnable_0;
  reg                 a_halted_fork2_logic_linkEnable_1;
  wire                when_Stream_l1094;
  wire                when_Stream_l1094_1;
  wire                a_cmdFork_fire;
  wire                a_dataFork_fire;
  reg        [1:0]    a_cmdFork_tracker_beat;
  wire                a_cmdFork_tracker_last;
  wire                when_Stream_l472;
  reg                 a_cmd_filtred_valid;
  wire                a_cmd_filtred_ready;
  wire       [2:0]    a_cmd_filtred_payload_opcode;
  wire       [2:0]    a_cmd_filtred_payload_param;
  wire       [1:0]    a_cmd_filtred_payload_source;
  wire       [31:0]   a_cmd_filtred_payload_address;
  wire       [2:0]    a_cmd_filtred_payload_size;
  wire       [15:0]   a_cmd_filtred_payload_mask;
  wire       [127:0]  a_cmd_filtred_payload_data;
  wire                a_cmd_filtred_payload_corrupt;
  wire                a_cmd_buffered_valid;
  wire                a_cmd_buffered_ready;
  wire       [2:0]    a_cmd_buffered_payload_opcode;
  wire       [2:0]    a_cmd_buffered_payload_param;
  wire       [1:0]    a_cmd_buffered_payload_source;
  wire       [31:0]   a_cmd_buffered_payload_address;
  wire       [2:0]    a_cmd_buffered_payload_size;
  wire       [15:0]   a_cmd_buffered_payload_mask;
  wire       [127:0]  a_cmd_buffered_payload_data;
  wire                a_cmd_buffered_payload_corrupt;
  reg                 a_cmd_filtred_rValid;
  wire                a_cmd_buffered_fire;
  reg        [2:0]    a_cmd_filtred_rData_opcode;
  reg        [2:0]    a_cmd_filtred_rData_param;
  reg        [1:0]    a_cmd_filtred_rData_source;
  reg        [31:0]   a_cmd_filtred_rData_address;
  reg        [2:0]    a_cmd_filtred_rData_size;
  reg        [15:0]   a_cmd_filtred_rData_mask;
  reg        [127:0]  a_cmd_filtred_rData_data;
  reg                 a_cmd_filtred_rData_corrupt;
  wire                a_cmd_isGet;
  wire       [7:0]    a_cmd_len;
  wire       [2:0]    a_cmd_sizePerBeat;
  wire                when_Stream_l472_1;
  reg                 a_data_filtred_valid;
  reg                 a_data_filtred_ready;
  wire       [2:0]    a_data_filtred_payload_opcode;
  wire       [2:0]    a_data_filtred_payload_param;
  wire       [1:0]    a_data_filtred_payload_source;
  wire       [31:0]   a_data_filtred_payload_address;
  wire       [2:0]    a_data_filtred_payload_size;
  wire       [15:0]   a_data_filtred_payload_mask;
  wire       [127:0]  a_data_filtred_payload_data;
  wire                a_data_filtred_payload_corrupt;
  wire                a_data_buffer_valid;
  wire                a_data_buffer_ready;
  wire       [2:0]    a_data_buffer_payload_opcode;
  wire       [2:0]    a_data_buffer_payload_param;
  wire       [1:0]    a_data_buffer_payload_source;
  wire       [31:0]   a_data_buffer_payload_address;
  wire       [2:0]    a_data_buffer_payload_size;
  wire       [15:0]   a_data_buffer_payload_mask;
  wire       [127:0]  a_data_buffer_payload_data;
  wire                a_data_buffer_payload_corrupt;
  reg                 a_data_filtred_rValid;
  reg        [2:0]    a_data_filtred_rData_opcode;
  reg        [2:0]    a_data_filtred_rData_param;
  reg        [1:0]    a_data_filtred_rData_source;
  reg        [31:0]   a_data_filtred_rData_address;
  reg        [2:0]    a_data_filtred_rData_size;
  reg        [15:0]   a_data_filtred_rData_mask;
  reg        [127:0]  a_data_filtred_rData_data;
  reg                 a_data_filtred_rData_corrupt;
  wire                when_Stream_l399;
  reg        [1:0]    a_data_buffer_tracker_beat;
  wire                a_data_buffer_tracker_last;
  wire                a_data_buffer_fire;
  wire       [2:0]    _zz_io_up_d_payload_opcode;
  `ifndef SYNTHESIS
  reg [127:0] io_up_a_payload_opcode_string;
  reg [119:0] io_up_d_payload_opcode_string;
  reg [127:0] a_halted_payload_opcode_string;
  reg [127:0] a_cmdFork_payload_opcode_string;
  reg [127:0] a_dataFork_payload_opcode_string;
  reg [127:0] a_cmd_filtred_payload_opcode_string;
  reg [127:0] a_cmd_buffered_payload_opcode_string;
  reg [127:0] a_cmd_filtred_rData_opcode_string;
  reg [127:0] a_data_filtred_payload_opcode_string;
  reg [127:0] a_data_buffer_payload_opcode_string;
  reg [127:0] a_data_filtred_rData_opcode_string;
  reg [119:0] _zz_io_up_d_payload_opcode_string;
  `endif


  ContextAsyncBufferFull a_ctx (
    .io_add_valid           (a_ctx_io_add_valid         ), //i
    .io_add_ready           (a_ctx_io_add_ready         ), //o
    .io_add_payload_id      (io_up_a_payload_source[1:0]), //i
    .io_add_payload_context (io_up_a_payload_size[2:0]  ), //i
    .io_remove_valid        (a_ctx_io_remove_valid      ), //i
    .io_remove_payload_id   (io_up_d_payload_source[1:0]), //i
    .io_query_id            (io_up_d_payload_source[1:0]), //i
    .io_query_context       (a_ctx_io_query_context[2:0]), //o
    .litex_clk              (litex_clk                  )  //i
  );
  StreamArbiter_7 d_arbiter (
    .io_inputs_0_valid          (io_down_b_valid                        ), //i
    .io_inputs_0_ready          (d_arbiter_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_source (io_down_b_payload_id[1:0]              ), //i
    .io_inputs_0_payload_denied (d_arbiter_io_inputs_0_payload_denied   ), //i
    .io_inputs_0_payload_last   (1'b1                                   ), //i
    .io_inputs_1_valid          (io_down_r_valid                        ), //i
    .io_inputs_1_ready          (d_arbiter_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_source (io_down_r_payload_id[1:0]              ), //i
    .io_inputs_1_payload_denied (d_arbiter_io_inputs_1_payload_denied   ), //i
    .io_inputs_1_payload_last   (io_down_r_payload_last                 ), //i
    .io_output_valid            (d_arbiter_io_output_valid              ), //o
    .io_output_ready            (io_up_d_ready                          ), //i
    .io_output_payload_source   (d_arbiter_io_output_payload_source[1:0]), //o
    .io_output_payload_denied   (d_arbiter_io_output_payload_denied     ), //o
    .io_output_payload_last     (d_arbiter_io_output_payload_last       ), //o
    .io_chosen                  (d_arbiter_io_chosen                    ), //o
    .io_chosenOH                (d_arbiter_io_chosenOH[1:0]             ), //o
    .litex_clk                  (litex_clk                              ), //i
    .cpuResetCtrl_reset         (cpuResetCtrl_reset                     )  //i
  );
  always @(*) begin
    case(io_up_a_payload_size)
      3'b000 : _zz_io_up_a_tracker_last = 2'b00;
      3'b001 : _zz_io_up_a_tracker_last = 2'b00;
      3'b010 : _zz_io_up_a_tracker_last = 2'b00;
      3'b011 : _zz_io_up_a_tracker_last = 2'b00;
      3'b100 : _zz_io_up_a_tracker_last = 2'b00;
      3'b101 : _zz_io_up_a_tracker_last = 2'b01;
      default : _zz_io_up_a_tracker_last = 2'b11;
    endcase
  end

  always @(*) begin
    case(io_up_d_payload_size)
      3'b000 : _zz_io_up_d_tracker_last = 2'b00;
      3'b001 : _zz_io_up_d_tracker_last = 2'b00;
      3'b010 : _zz_io_up_d_tracker_last = 2'b00;
      3'b011 : _zz_io_up_d_tracker_last = 2'b00;
      3'b100 : _zz_io_up_d_tracker_last = 2'b00;
      3'b101 : _zz_io_up_d_tracker_last = 2'b01;
      default : _zz_io_up_d_tracker_last = 2'b11;
    endcase
  end

  always @(*) begin
    case(a_cmdFork_payload_size)
      3'b000 : _zz_a_cmdFork_tracker_last = 2'b00;
      3'b001 : _zz_a_cmdFork_tracker_last = 2'b00;
      3'b010 : _zz_a_cmdFork_tracker_last = 2'b00;
      3'b011 : _zz_a_cmdFork_tracker_last = 2'b00;
      3'b100 : _zz_a_cmdFork_tracker_last = 2'b00;
      3'b101 : _zz_a_cmdFork_tracker_last = 2'b01;
      default : _zz_a_cmdFork_tracker_last = 2'b11;
    endcase
  end

  always @(*) begin
    case(a_cmd_buffered_payload_size)
      3'b000 : begin
        _zz_a_cmd_len = 2'b00;
        _zz_a_cmd_sizePerBeat = 3'b000;
      end
      3'b001 : begin
        _zz_a_cmd_len = 2'b00;
        _zz_a_cmd_sizePerBeat = 3'b001;
      end
      3'b010 : begin
        _zz_a_cmd_len = 2'b00;
        _zz_a_cmd_sizePerBeat = 3'b010;
      end
      3'b011 : begin
        _zz_a_cmd_len = 2'b00;
        _zz_a_cmd_sizePerBeat = 3'b011;
      end
      3'b100 : begin
        _zz_a_cmd_len = 2'b00;
        _zz_a_cmd_sizePerBeat = 3'b100;
      end
      3'b101 : begin
        _zz_a_cmd_len = 2'b01;
        _zz_a_cmd_sizePerBeat = 3'b100;
      end
      default : begin
        _zz_a_cmd_len = 2'b11;
        _zz_a_cmd_sizePerBeat = 3'b100;
      end
    endcase
  end

  always @(*) begin
    case(a_data_buffer_payload_size)
      3'b000 : _zz_a_data_buffer_tracker_last = 2'b00;
      3'b001 : _zz_a_data_buffer_tracker_last = 2'b00;
      3'b010 : _zz_a_data_buffer_tracker_last = 2'b00;
      3'b011 : _zz_a_data_buffer_tracker_last = 2'b00;
      3'b100 : _zz_a_data_buffer_tracker_last = 2'b00;
      3'b101 : _zz_a_data_buffer_tracker_last = 2'b01;
      default : _zz_a_data_buffer_tracker_last = 2'b11;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_up_a_payload_opcode)
      A_PUT_FULL_DATA : io_up_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_up_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_up_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_up_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_up_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_up_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_up_d_payload_opcode)
      D_ACCESS_ACK : io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(a_halted_payload_opcode)
      A_PUT_FULL_DATA : a_halted_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_halted_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_halted_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_halted_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_halted_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_halted_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmdFork_payload_opcode)
      A_PUT_FULL_DATA : a_cmdFork_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmdFork_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmdFork_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmdFork_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmdFork_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmdFork_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_dataFork_payload_opcode)
      A_PUT_FULL_DATA : a_dataFork_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_dataFork_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_dataFork_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_dataFork_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_dataFork_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_dataFork_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmd_filtred_payload_opcode)
      A_PUT_FULL_DATA : a_cmd_filtred_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmd_filtred_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmd_filtred_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmd_filtred_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmd_filtred_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmd_filtred_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmd_buffered_payload_opcode)
      A_PUT_FULL_DATA : a_cmd_buffered_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmd_buffered_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmd_buffered_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmd_buffered_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmd_buffered_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmd_buffered_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_cmd_filtred_rData_opcode)
      A_PUT_FULL_DATA : a_cmd_filtred_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_cmd_filtred_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_cmd_filtred_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_cmd_filtred_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_cmd_filtred_rData_opcode_string = "ACQUIRE_PERM    ";
      default : a_cmd_filtred_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_data_filtred_payload_opcode)
      A_PUT_FULL_DATA : a_data_filtred_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_data_filtred_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_data_filtred_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_data_filtred_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_data_filtred_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_data_filtred_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_data_buffer_payload_opcode)
      A_PUT_FULL_DATA : a_data_buffer_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_data_buffer_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_data_buffer_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_data_buffer_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_data_buffer_payload_opcode_string = "ACQUIRE_PERM    ";
      default : a_data_buffer_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(a_data_filtred_rData_opcode)
      A_PUT_FULL_DATA : a_data_filtred_rData_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : a_data_filtred_rData_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : a_data_filtred_rData_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : a_data_filtred_rData_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : a_data_filtred_rData_opcode_string = "ACQUIRE_PERM    ";
      default : a_data_filtred_rData_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_up_d_payload_opcode)
      D_ACCESS_ACK : _zz_io_up_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_up_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_up_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_up_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_up_d_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_up_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  always @(*) begin
    a_ctxFull = 1'b0;
    if(when_ContextBuffer_l19) begin
      a_ctxFull = 1'b1;
    end
  end

  assign _zz_io_up_a_ready = (! a_ctxFull);
  assign a_halted_valid = (io_up_a_valid && _zz_io_up_a_ready);
  assign io_up_a_ready = (a_halted_ready && _zz_io_up_a_ready);
  assign a_halted_payload_opcode = io_up_a_payload_opcode;
  assign a_halted_payload_param = io_up_a_payload_param;
  assign a_halted_payload_source = io_up_a_payload_source;
  assign a_halted_payload_address = io_up_a_payload_address;
  assign a_halted_payload_size = io_up_a_payload_size;
  assign a_halted_payload_mask = io_up_a_payload_mask;
  assign a_halted_payload_data = io_up_a_payload_data;
  assign a_halted_payload_corrupt = io_up_a_payload_corrupt;
  assign io_up_a_fire = (io_up_a_valid && io_up_a_ready);
  assign io_up_a_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == io_up_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_up_a_payload_opcode))) || (io_up_a_tracker_beat == _zz_io_up_a_tracker_last));
  assign a_ctx_io_add_valid = (io_up_a_fire && io_up_a_tracker_last);
  assign when_ContextBuffer_l19 = (! a_ctx_io_add_ready);
  assign io_up_d_fire = (io_up_d_valid && io_up_d_ready);
  assign io_up_d_tracker_last = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_up_d_payload_opcode)) || (D_GRANT_DATA == io_up_d_payload_opcode))) || (io_up_d_tracker_beat == _zz_io_up_d_tracker_last));
  assign a_ctx_io_remove_valid = ((io_up_d_fire && io_up_d_tracker_last) && (|{(io_up_d_payload_opcode == D_GRANT_DATA),{(io_up_d_payload_opcode == D_GRANT),{(io_up_d_payload_opcode == D_ACCESS_ACK_DATA),(io_up_d_payload_opcode == D_ACCESS_ACK)}}}));
  always @(*) begin
    a_halted_ready = 1'b1;
    if(when_Stream_l1094) begin
      a_halted_ready = 1'b0;
    end
    if(when_Stream_l1094_1) begin
      a_halted_ready = 1'b0;
    end
  end

  assign when_Stream_l1094 = ((! a_cmdFork_ready) && a_halted_fork2_logic_linkEnable_0);
  assign when_Stream_l1094_1 = ((! a_dataFork_ready) && a_halted_fork2_logic_linkEnable_1);
  assign a_cmdFork_valid = (a_halted_valid && a_halted_fork2_logic_linkEnable_0);
  assign a_cmdFork_payload_opcode = a_halted_payload_opcode;
  assign a_cmdFork_payload_param = a_halted_payload_param;
  assign a_cmdFork_payload_source = a_halted_payload_source;
  assign a_cmdFork_payload_address = a_halted_payload_address;
  assign a_cmdFork_payload_size = a_halted_payload_size;
  assign a_cmdFork_payload_mask = a_halted_payload_mask;
  assign a_cmdFork_payload_data = a_halted_payload_data;
  assign a_cmdFork_payload_corrupt = a_halted_payload_corrupt;
  assign a_cmdFork_fire = (a_cmdFork_valid && a_cmdFork_ready);
  assign a_dataFork_valid = (a_halted_valid && a_halted_fork2_logic_linkEnable_1);
  assign a_dataFork_payload_opcode = a_halted_payload_opcode;
  assign a_dataFork_payload_param = a_halted_payload_param;
  assign a_dataFork_payload_source = a_halted_payload_source;
  assign a_dataFork_payload_address = a_halted_payload_address;
  assign a_dataFork_payload_size = a_halted_payload_size;
  assign a_dataFork_payload_mask = a_halted_payload_mask;
  assign a_dataFork_payload_data = a_halted_payload_data;
  assign a_dataFork_payload_corrupt = a_halted_payload_corrupt;
  assign a_dataFork_fire = (a_dataFork_valid && a_dataFork_ready);
  assign a_cmdFork_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == a_cmdFork_payload_opcode)) || (A_PUT_PARTIAL_DATA == a_cmdFork_payload_opcode))) || (a_cmdFork_tracker_beat == _zz_a_cmdFork_tracker_last));
  assign when_Stream_l472 = (! (a_cmdFork_tracker_beat == 2'b00));
  always @(*) begin
    a_cmd_filtred_valid = a_cmdFork_valid;
    if(when_Stream_l472) begin
      a_cmd_filtred_valid = 1'b0;
    end
  end

  always @(*) begin
    a_cmdFork_ready = a_cmd_filtred_ready;
    if(when_Stream_l472) begin
      a_cmdFork_ready = 1'b1;
    end
  end

  assign a_cmd_filtred_payload_opcode = a_cmdFork_payload_opcode;
  assign a_cmd_filtred_payload_param = a_cmdFork_payload_param;
  assign a_cmd_filtred_payload_source = a_cmdFork_payload_source;
  assign a_cmd_filtred_payload_address = a_cmdFork_payload_address;
  assign a_cmd_filtred_payload_size = a_cmdFork_payload_size;
  assign a_cmd_filtred_payload_mask = a_cmdFork_payload_mask;
  assign a_cmd_filtred_payload_data = a_cmdFork_payload_data;
  assign a_cmd_filtred_payload_corrupt = a_cmdFork_payload_corrupt;
  assign a_cmd_buffered_fire = (a_cmd_buffered_valid && a_cmd_buffered_ready);
  assign a_cmd_filtred_ready = (! a_cmd_filtred_rValid);
  assign a_cmd_buffered_valid = a_cmd_filtred_rValid;
  assign a_cmd_buffered_payload_opcode = a_cmd_filtred_rData_opcode;
  assign a_cmd_buffered_payload_param = a_cmd_filtred_rData_param;
  assign a_cmd_buffered_payload_source = a_cmd_filtred_rData_source;
  assign a_cmd_buffered_payload_address = a_cmd_filtred_rData_address;
  assign a_cmd_buffered_payload_size = a_cmd_filtred_rData_size;
  assign a_cmd_buffered_payload_mask = a_cmd_filtred_rData_mask;
  assign a_cmd_buffered_payload_data = a_cmd_filtred_rData_data;
  assign a_cmd_buffered_payload_corrupt = a_cmd_filtred_rData_corrupt;
  assign a_cmd_isGet = (a_cmd_buffered_payload_opcode == A_GET);
  assign io_down_aw_valid = (a_cmd_buffered_valid && (! a_cmd_isGet));
  assign io_down_ar_valid = (a_cmd_buffered_valid && a_cmd_isGet);
  assign a_cmd_buffered_ready = (a_cmd_isGet ? io_down_ar_ready : io_down_aw_ready);
  assign a_cmd_len = {6'd0, _zz_a_cmd_len};
  assign a_cmd_sizePerBeat = _zz_a_cmd_sizePerBeat;
  assign io_down_aw_payload_addr = a_cmd_buffered_payload_address;
  assign io_down_aw_payload_id = a_cmd_buffered_payload_source;
  assign io_down_aw_payload_len = a_cmd_len;
  assign io_down_aw_payload_size = a_cmd_sizePerBeat;
  assign io_down_aw_payload_burst = 2'b01;
  assign io_down_ar_payload_addr = a_cmd_buffered_payload_address;
  assign io_down_ar_payload_id = a_cmd_buffered_payload_source;
  assign io_down_ar_payload_len = a_cmd_len;
  assign io_down_ar_payload_size = a_cmd_sizePerBeat;
  assign io_down_ar_payload_burst = 2'b01;
  assign io_down_aw_payload_allStrb = (a_cmd_buffered_payload_opcode == A_PUT_FULL_DATA);
  assign when_Stream_l472_1 = (! ((a_dataFork_payload_opcode == A_PUT_FULL_DATA) || (a_dataFork_payload_opcode == A_PUT_PARTIAL_DATA)));
  always @(*) begin
    a_data_filtred_valid = a_dataFork_valid;
    if(when_Stream_l472_1) begin
      a_data_filtred_valid = 1'b0;
    end
  end

  always @(*) begin
    a_dataFork_ready = a_data_filtred_ready;
    if(when_Stream_l472_1) begin
      a_dataFork_ready = 1'b1;
    end
  end

  assign a_data_filtred_payload_opcode = a_dataFork_payload_opcode;
  assign a_data_filtred_payload_param = a_dataFork_payload_param;
  assign a_data_filtred_payload_source = a_dataFork_payload_source;
  assign a_data_filtred_payload_address = a_dataFork_payload_address;
  assign a_data_filtred_payload_size = a_dataFork_payload_size;
  assign a_data_filtred_payload_mask = a_dataFork_payload_mask;
  assign a_data_filtred_payload_data = a_dataFork_payload_data;
  assign a_data_filtred_payload_corrupt = a_dataFork_payload_corrupt;
  always @(*) begin
    a_data_filtred_ready = a_data_buffer_ready;
    if(when_Stream_l399) begin
      a_data_filtred_ready = 1'b1;
    end
  end

  assign when_Stream_l399 = (! a_data_buffer_valid);
  assign a_data_buffer_valid = a_data_filtred_rValid;
  assign a_data_buffer_payload_opcode = a_data_filtred_rData_opcode;
  assign a_data_buffer_payload_param = a_data_filtred_rData_param;
  assign a_data_buffer_payload_source = a_data_filtred_rData_source;
  assign a_data_buffer_payload_address = a_data_filtred_rData_address;
  assign a_data_buffer_payload_size = a_data_filtred_rData_size;
  assign a_data_buffer_payload_mask = a_data_filtred_rData_mask;
  assign a_data_buffer_payload_data = a_data_filtred_rData_data;
  assign a_data_buffer_payload_corrupt = a_data_filtred_rData_corrupt;
  assign io_down_w_valid = a_data_buffer_valid;
  assign a_data_buffer_ready = io_down_w_ready;
  assign io_down_w_payload_data = a_data_buffer_payload_data;
  assign io_down_w_payload_strb = a_data_buffer_payload_mask;
  assign a_data_buffer_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == a_data_buffer_payload_opcode)) || (A_PUT_PARTIAL_DATA == a_data_buffer_payload_opcode))) || (a_data_buffer_tracker_beat == _zz_a_data_buffer_tracker_last));
  assign a_data_buffer_fire = (a_data_buffer_valid && a_data_buffer_ready);
  assign io_down_w_payload_last = a_data_buffer_tracker_last;
  assign io_down_b_ready = d_arbiter_io_inputs_0_ready;
  assign d_arbiter_io_inputs_0_payload_denied = (! (io_down_b_payload_resp == 2'b00));
  assign io_down_r_ready = d_arbiter_io_inputs_1_ready;
  assign d_arbiter_io_inputs_1_payload_denied = (! (io_down_r_payload_resp == 2'b00));
  assign io_up_d_valid = d_arbiter_io_output_valid;
  assign _zz_io_up_d_payload_opcode = (d_arbiter_io_chosen[0] ? D_ACCESS_ACK_DATA : D_ACCESS_ACK);
  assign io_up_d_payload_opcode = _zz_io_up_d_payload_opcode;
  assign io_up_d_payload_param = 3'b000;
  assign io_up_d_payload_source = d_arbiter_io_output_payload_source;
  assign io_up_d_payload_denied = d_arbiter_io_output_payload_denied;
  assign io_up_d_payload_data = io_down_r_payload_data;
  assign io_up_d_payload_corrupt = 1'b0;
  assign io_up_d_payload_size = a_ctx_io_query_context;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      io_up_a_tracker_beat <= 2'b00;
      io_up_d_tracker_beat <= 2'b00;
      a_halted_fork2_logic_linkEnable_0 <= 1'b1;
      a_halted_fork2_logic_linkEnable_1 <= 1'b1;
      a_cmdFork_tracker_beat <= 2'b00;
      a_cmd_filtred_rValid <= 1'b0;
      a_data_filtred_rValid <= 1'b0;
      a_data_buffer_tracker_beat <= 2'b00;
    end else begin
      if(io_up_a_fire) begin
        io_up_a_tracker_beat <= (io_up_a_tracker_beat + 2'b01);
        if(io_up_a_tracker_last) begin
          io_up_a_tracker_beat <= 2'b00;
        end
      end
      if(io_up_d_fire) begin
        io_up_d_tracker_beat <= (io_up_d_tracker_beat + 2'b01);
        if(io_up_d_tracker_last) begin
          io_up_d_tracker_beat <= 2'b00;
        end
      end
      if(a_cmdFork_fire) begin
        a_halted_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(a_dataFork_fire) begin
        a_halted_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(a_halted_ready) begin
        a_halted_fork2_logic_linkEnable_0 <= 1'b1;
        a_halted_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(a_cmdFork_fire) begin
        a_cmdFork_tracker_beat <= (a_cmdFork_tracker_beat + 2'b01);
        if(a_cmdFork_tracker_last) begin
          a_cmdFork_tracker_beat <= 2'b00;
        end
      end
      if(a_cmd_filtred_valid) begin
        a_cmd_filtred_rValid <= 1'b1;
      end
      if(a_cmd_buffered_fire) begin
        a_cmd_filtred_rValid <= 1'b0;
      end
      if(a_data_filtred_ready) begin
        a_data_filtred_rValid <= a_data_filtred_valid;
      end
      if(a_data_buffer_fire) begin
        a_data_buffer_tracker_beat <= (a_data_buffer_tracker_beat + 2'b01);
        if(a_data_buffer_tracker_last) begin
          a_data_buffer_tracker_beat <= 2'b00;
        end
      end
    end
  end

  always @(posedge litex_clk) begin
    if(a_cmd_filtred_ready) begin
      a_cmd_filtred_rData_opcode <= a_cmd_filtred_payload_opcode;
      a_cmd_filtred_rData_param <= a_cmd_filtred_payload_param;
      a_cmd_filtred_rData_source <= a_cmd_filtred_payload_source;
      a_cmd_filtred_rData_address <= a_cmd_filtred_payload_address;
      a_cmd_filtred_rData_size <= a_cmd_filtred_payload_size;
      a_cmd_filtred_rData_mask <= a_cmd_filtred_payload_mask;
      a_cmd_filtred_rData_data <= a_cmd_filtred_payload_data;
      a_cmd_filtred_rData_corrupt <= a_cmd_filtred_payload_corrupt;
    end
    if(a_data_filtred_ready) begin
      a_data_filtred_rData_opcode <= a_data_filtred_payload_opcode;
      a_data_filtred_rData_param <= a_data_filtred_payload_param;
      a_data_filtred_rData_source <= a_data_filtred_payload_source;
      a_data_filtred_rData_address <= a_data_filtred_payload_address;
      a_data_filtred_rData_size <= a_data_filtred_payload_size;
      a_data_filtred_rData_mask <= a_data_filtred_payload_mask;
      a_data_filtred_rData_data <= a_data_filtred_payload_data;
      a_data_filtred_rData_corrupt <= a_data_filtred_payload_corrupt;
    end
  end


endmodule

module Arbiter_1 (
  input  wire          io_ups_0_a_valid,
  output wire          io_ups_0_a_ready,
  input  wire [2:0]    io_ups_0_a_payload_opcode,
  input  wire [2:0]    io_ups_0_a_payload_param,
  input  wire [31:0]   io_ups_0_a_payload_address,
  input  wire [1:0]    io_ups_0_a_payload_size,
  input  wire [3:0]    io_ups_0_a_payload_mask,
  input  wire [31:0]   io_ups_0_a_payload_data,
  input  wire          io_ups_0_a_payload_corrupt,
  output wire          io_ups_0_d_valid,
  input  wire          io_ups_0_d_ready,
  output wire [2:0]    io_ups_0_d_payload_opcode,
  output wire [2:0]    io_ups_0_d_payload_param,
  output wire [1:0]    io_ups_0_d_payload_size,
  output wire          io_ups_0_d_payload_denied,
  output wire [31:0]   io_ups_0_d_payload_data,
  output wire          io_ups_0_d_payload_corrupt,
  input  wire          io_ups_1_a_valid,
  output wire          io_ups_1_a_ready,
  input  wire [2:0]    io_ups_1_a_payload_opcode,
  input  wire [2:0]    io_ups_1_a_payload_param,
  input  wire [1:0]    io_ups_1_a_payload_source,
  input  wire [31:0]   io_ups_1_a_payload_address,
  input  wire [2:0]    io_ups_1_a_payload_size,
  input  wire [3:0]    io_ups_1_a_payload_mask,
  input  wire [31:0]   io_ups_1_a_payload_data,
  input  wire          io_ups_1_a_payload_corrupt,
  output wire          io_ups_1_d_valid,
  input  wire          io_ups_1_d_ready,
  output wire [2:0]    io_ups_1_d_payload_opcode,
  output wire [2:0]    io_ups_1_d_payload_param,
  output wire [1:0]    io_ups_1_d_payload_source,
  output wire [2:0]    io_ups_1_d_payload_size,
  output wire          io_ups_1_d_payload_denied,
  output wire [31:0]   io_ups_1_d_payload_data,
  output wire          io_ups_1_d_payload_corrupt,
  output wire          io_down_a_valid,
  input  wire          io_down_a_ready,
  output wire [2:0]    io_down_a_payload_opcode,
  output wire [2:0]    io_down_a_payload_param,
  output wire [2:0]    io_down_a_payload_source,
  output wire [31:0]   io_down_a_payload_address,
  output wire [2:0]    io_down_a_payload_size,
  output wire [3:0]    io_down_a_payload_mask,
  output wire [31:0]   io_down_a_payload_data,
  output wire          io_down_a_payload_corrupt,
  input  wire          io_down_d_valid,
  output wire          io_down_d_ready,
  input  wire [2:0]    io_down_d_payload_opcode,
  input  wire [2:0]    io_down_d_payload_param,
  input  wire [2:0]    io_down_d_payload_source,
  input  wire [2:0]    io_down_d_payload_size,
  input  wire          io_down_d_payload_denied,
  input  wire [31:0]   io_down_d_payload_data,
  input  wire          io_down_d_payload_corrupt,
  input  wire          litex_clk,
  input  wire          litex_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire       [2:0]    a_arbiter_io_inputs_0_payload_size;
  wire                a_arbiter_io_inputs_0_ready;
  wire                a_arbiter_io_inputs_1_ready;
  wire                a_arbiter_io_output_valid;
  wire       [2:0]    a_arbiter_io_output_payload_opcode;
  wire       [2:0]    a_arbiter_io_output_payload_param;
  wire       [2:0]    a_arbiter_io_output_payload_source;
  wire       [31:0]   a_arbiter_io_output_payload_address;
  wire       [2:0]    a_arbiter_io_output_payload_size;
  wire       [3:0]    a_arbiter_io_output_payload_mask;
  wire       [31:0]   a_arbiter_io_output_payload_data;
  wire                a_arbiter_io_output_payload_corrupt;
  wire       [0:0]    a_arbiter_io_chosen;
  wire       [1:0]    a_arbiter_io_chosenOH;
  wire       [2:0]    _zz_ups_1_a_payload_source;
  reg                 _zz_io_down_d_ready;
  wire                ups_0_a_valid;
  wire                ups_0_a_ready;
  wire       [2:0]    ups_0_a_payload_opcode;
  wire       [2:0]    ups_0_a_payload_param;
  wire       [2:0]    ups_0_a_payload_source;
  wire       [31:0]   ups_0_a_payload_address;
  wire       [1:0]    ups_0_a_payload_size;
  wire       [3:0]    ups_0_a_payload_mask;
  wire       [31:0]   ups_0_a_payload_data;
  wire                ups_0_a_payload_corrupt;
  wire                ups_0_d_valid;
  wire                ups_0_d_ready;
  wire       [2:0]    ups_0_d_payload_opcode;
  wire       [2:0]    ups_0_d_payload_param;
  wire       [2:0]    ups_0_d_payload_source;
  wire       [1:0]    ups_0_d_payload_size;
  wire                ups_0_d_payload_denied;
  wire       [31:0]   ups_0_d_payload_data;
  wire                ups_0_d_payload_corrupt;
  wire                ups_1_a_valid;
  wire                ups_1_a_ready;
  wire       [2:0]    ups_1_a_payload_opcode;
  wire       [2:0]    ups_1_a_payload_param;
  wire       [2:0]    ups_1_a_payload_source;
  wire       [31:0]   ups_1_a_payload_address;
  wire       [2:0]    ups_1_a_payload_size;
  wire       [3:0]    ups_1_a_payload_mask;
  wire       [31:0]   ups_1_a_payload_data;
  wire                ups_1_a_payload_corrupt;
  wire                ups_1_d_valid;
  wire                ups_1_d_ready;
  wire       [2:0]    ups_1_d_payload_opcode;
  wire       [2:0]    ups_1_d_payload_param;
  wire       [2:0]    ups_1_d_payload_source;
  wire       [2:0]    ups_1_d_payload_size;
  wire                ups_1_d_payload_denied;
  wire       [31:0]   ups_1_d_payload_data;
  wire                ups_1_d_payload_corrupt;
  wire       [0:0]    d_sel;
  `ifndef SYNTHESIS
  reg [127:0] io_ups_0_a_payload_opcode_string;
  reg [119:0] io_ups_0_d_payload_opcode_string;
  reg [127:0] io_ups_1_a_payload_opcode_string;
  reg [119:0] io_ups_1_d_payload_opcode_string;
  reg [127:0] io_down_a_payload_opcode_string;
  reg [119:0] io_down_d_payload_opcode_string;
  reg [127:0] ups_0_a_payload_opcode_string;
  reg [119:0] ups_0_d_payload_opcode_string;
  reg [127:0] ups_1_a_payload_opcode_string;
  reg [119:0] ups_1_d_payload_opcode_string;
  `endif


  assign _zz_ups_1_a_payload_source = {1'd0, io_ups_1_a_payload_source};
  StreamArbiter_6 a_arbiter (
    .io_inputs_0_valid           (ups_0_a_valid                            ), //i
    .io_inputs_0_ready           (a_arbiter_io_inputs_0_ready              ), //o
    .io_inputs_0_payload_opcode  (ups_0_a_payload_opcode[2:0]              ), //i
    .io_inputs_0_payload_param   (ups_0_a_payload_param[2:0]               ), //i
    .io_inputs_0_payload_source  (ups_0_a_payload_source[2:0]              ), //i
    .io_inputs_0_payload_address (ups_0_a_payload_address[31:0]            ), //i
    .io_inputs_0_payload_size    (a_arbiter_io_inputs_0_payload_size[2:0]  ), //i
    .io_inputs_0_payload_mask    (ups_0_a_payload_mask[3:0]                ), //i
    .io_inputs_0_payload_data    (ups_0_a_payload_data[31:0]               ), //i
    .io_inputs_0_payload_corrupt (ups_0_a_payload_corrupt                  ), //i
    .io_inputs_1_valid           (ups_1_a_valid                            ), //i
    .io_inputs_1_ready           (a_arbiter_io_inputs_1_ready              ), //o
    .io_inputs_1_payload_opcode  (ups_1_a_payload_opcode[2:0]              ), //i
    .io_inputs_1_payload_param   (ups_1_a_payload_param[2:0]               ), //i
    .io_inputs_1_payload_source  (ups_1_a_payload_source[2:0]              ), //i
    .io_inputs_1_payload_address (ups_1_a_payload_address[31:0]            ), //i
    .io_inputs_1_payload_size    (ups_1_a_payload_size[2:0]                ), //i
    .io_inputs_1_payload_mask    (ups_1_a_payload_mask[3:0]                ), //i
    .io_inputs_1_payload_data    (ups_1_a_payload_data[31:0]               ), //i
    .io_inputs_1_payload_corrupt (ups_1_a_payload_corrupt                  ), //i
    .io_output_valid             (a_arbiter_io_output_valid                ), //o
    .io_output_ready             (io_down_a_ready                          ), //i
    .io_output_payload_opcode    (a_arbiter_io_output_payload_opcode[2:0]  ), //o
    .io_output_payload_param     (a_arbiter_io_output_payload_param[2:0]   ), //o
    .io_output_payload_source    (a_arbiter_io_output_payload_source[2:0]  ), //o
    .io_output_payload_address   (a_arbiter_io_output_payload_address[31:0]), //o
    .io_output_payload_size      (a_arbiter_io_output_payload_size[2:0]    ), //o
    .io_output_payload_mask      (a_arbiter_io_output_payload_mask[3:0]    ), //o
    .io_output_payload_data      (a_arbiter_io_output_payload_data[31:0]   ), //o
    .io_output_payload_corrupt   (a_arbiter_io_output_payload_corrupt      ), //o
    .io_chosen                   (a_arbiter_io_chosen                      ), //o
    .io_chosenOH                 (a_arbiter_io_chosenOH[1:0]               ), //o
    .litex_clk                   (litex_clk                                ), //i
    .litex_reset                 (litex_reset                              )  //i
  );
  always @(*) begin
    case(d_sel)
      1'b0 : _zz_io_down_d_ready = ups_0_d_ready;
      default : _zz_io_down_d_ready = ups_1_d_ready;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_ups_0_a_payload_opcode)
      A_PUT_FULL_DATA : io_ups_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_ups_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_ups_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_ups_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_ups_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_ups_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_0_d_payload_opcode)
      D_ACCESS_ACK : io_ups_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_ups_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_ups_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_ups_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_ups_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_ups_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_1_a_payload_opcode)
      A_PUT_FULL_DATA : io_ups_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_ups_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_ups_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_ups_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_ups_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_ups_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_1_d_payload_opcode)
      D_ACCESS_ACK : io_ups_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_ups_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_ups_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_ups_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_ups_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_ups_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_down_a_payload_opcode)
      A_PUT_FULL_DATA : io_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_down_d_payload_opcode)
      D_ACCESS_ACK : io_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ups_0_a_payload_opcode)
      A_PUT_FULL_DATA : ups_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ups_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ups_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ups_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ups_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ups_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ups_0_d_payload_opcode)
      D_ACCESS_ACK : ups_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ups_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ups_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ups_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ups_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ups_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ups_1_a_payload_opcode)
      A_PUT_FULL_DATA : ups_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ups_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ups_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ups_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ups_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ups_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ups_1_d_payload_opcode)
      D_ACCESS_ACK : ups_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ups_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ups_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ups_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ups_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ups_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign ups_0_a_valid = io_ups_0_a_valid;
  assign io_ups_0_a_ready = ups_0_a_ready;
  assign ups_0_a_payload_opcode = io_ups_0_a_payload_opcode;
  assign ups_0_a_payload_param = io_ups_0_a_payload_param;
  assign ups_0_a_payload_address = io_ups_0_a_payload_address;
  assign ups_0_a_payload_size = io_ups_0_a_payload_size;
  assign ups_0_a_payload_mask = io_ups_0_a_payload_mask;
  assign ups_0_a_payload_data = io_ups_0_a_payload_data;
  assign ups_0_a_payload_corrupt = io_ups_0_a_payload_corrupt;
  assign io_ups_0_d_valid = ups_0_d_valid;
  assign ups_0_d_ready = io_ups_0_d_ready;
  assign io_ups_0_d_payload_opcode = ups_0_d_payload_opcode;
  assign io_ups_0_d_payload_param = ups_0_d_payload_param;
  assign io_ups_0_d_payload_size = ups_0_d_payload_size;
  assign io_ups_0_d_payload_denied = ups_0_d_payload_denied;
  assign io_ups_0_d_payload_data = ups_0_d_payload_data;
  assign io_ups_0_d_payload_corrupt = ups_0_d_payload_corrupt;
  assign ups_0_a_payload_source = (3'b000 | 3'b000);
  assign ups_1_a_valid = io_ups_1_a_valid;
  assign io_ups_1_a_ready = ups_1_a_ready;
  assign ups_1_a_payload_opcode = io_ups_1_a_payload_opcode;
  assign ups_1_a_payload_param = io_ups_1_a_payload_param;
  assign ups_1_a_payload_address = io_ups_1_a_payload_address;
  assign ups_1_a_payload_size = io_ups_1_a_payload_size;
  assign ups_1_a_payload_mask = io_ups_1_a_payload_mask;
  assign ups_1_a_payload_data = io_ups_1_a_payload_data;
  assign ups_1_a_payload_corrupt = io_ups_1_a_payload_corrupt;
  assign io_ups_1_d_valid = ups_1_d_valid;
  assign ups_1_d_ready = io_ups_1_d_ready;
  assign io_ups_1_d_payload_opcode = ups_1_d_payload_opcode;
  assign io_ups_1_d_payload_param = ups_1_d_payload_param;
  assign io_ups_1_d_payload_size = ups_1_d_payload_size;
  assign io_ups_1_d_payload_denied = ups_1_d_payload_denied;
  assign io_ups_1_d_payload_data = ups_1_d_payload_data;
  assign io_ups_1_d_payload_corrupt = ups_1_d_payload_corrupt;
  assign ups_1_a_payload_source = (_zz_ups_1_a_payload_source | 3'b100);
  assign io_ups_1_d_payload_source = ups_1_d_payload_source[1:0];
  assign ups_0_a_ready = a_arbiter_io_inputs_0_ready;
  assign a_arbiter_io_inputs_0_payload_size = {1'd0, ups_0_a_payload_size};
  assign ups_1_a_ready = a_arbiter_io_inputs_1_ready;
  assign io_down_a_valid = a_arbiter_io_output_valid;
  assign io_down_a_payload_opcode = a_arbiter_io_output_payload_opcode;
  assign io_down_a_payload_param = a_arbiter_io_output_payload_param;
  assign io_down_a_payload_source = a_arbiter_io_output_payload_source;
  assign io_down_a_payload_address = a_arbiter_io_output_payload_address;
  assign io_down_a_payload_size = a_arbiter_io_output_payload_size;
  assign io_down_a_payload_mask = a_arbiter_io_output_payload_mask;
  assign io_down_a_payload_data = a_arbiter_io_output_payload_data;
  assign io_down_a_payload_corrupt = a_arbiter_io_output_payload_corrupt;
  assign d_sel = io_down_d_payload_source[2 : 2];
  assign io_down_d_ready = _zz_io_down_d_ready;
  assign ups_0_d_valid = (io_down_d_valid && (d_sel == 1'b0));
  assign ups_0_d_payload_opcode = io_down_d_payload_opcode;
  assign ups_0_d_payload_param = io_down_d_payload_param;
  assign ups_0_d_payload_source = io_down_d_payload_source;
  assign ups_0_d_payload_denied = io_down_d_payload_denied;
  assign ups_0_d_payload_size = io_down_d_payload_size[1:0];
  assign ups_0_d_payload_data = io_down_d_payload_data;
  assign ups_0_d_payload_corrupt = io_down_d_payload_corrupt;
  assign ups_1_d_valid = (io_down_d_valid && (d_sel == 1'b1));
  assign ups_1_d_payload_opcode = io_down_d_payload_opcode;
  assign ups_1_d_payload_param = io_down_d_payload_param;
  assign ups_1_d_payload_source = io_down_d_payload_source;
  assign ups_1_d_payload_denied = io_down_d_payload_denied;
  assign ups_1_d_payload_size = io_down_d_payload_size;
  assign ups_1_d_payload_data = io_down_d_payload_data;
  assign ups_1_d_payload_corrupt = io_down_d_payload_corrupt;

endmodule

module Arbiter (
  input  wire          io_ups_0_a_valid,
  output wire          io_ups_0_a_ready,
  input  wire [2:0]    io_ups_0_a_payload_opcode,
  input  wire [2:0]    io_ups_0_a_payload_param,
  input  wire [31:0]   io_ups_0_a_payload_address,
  input  wire [2:0]    io_ups_0_a_payload_size,
  output wire          io_ups_0_d_valid,
  input  wire          io_ups_0_d_ready,
  output wire [2:0]    io_ups_0_d_payload_opcode,
  output wire [2:0]    io_ups_0_d_payload_param,
  output wire [2:0]    io_ups_0_d_payload_size,
  output wire          io_ups_0_d_payload_denied,
  output wire [63:0]   io_ups_0_d_payload_data,
  output wire          io_ups_0_d_payload_corrupt,
  input  wire          io_ups_1_a_valid,
  output wire          io_ups_1_a_ready,
  input  wire [2:0]    io_ups_1_a_payload_opcode,
  input  wire [2:0]    io_ups_1_a_payload_param,
  input  wire [0:0]    io_ups_1_a_payload_source,
  input  wire [31:0]   io_ups_1_a_payload_address,
  input  wire [2:0]    io_ups_1_a_payload_size,
  input  wire [7:0]    io_ups_1_a_payload_mask,
  input  wire [63:0]   io_ups_1_a_payload_data,
  input  wire          io_ups_1_a_payload_corrupt,
  output wire          io_ups_1_d_valid,
  input  wire          io_ups_1_d_ready,
  output wire [2:0]    io_ups_1_d_payload_opcode,
  output wire [2:0]    io_ups_1_d_payload_param,
  output wire [0:0]    io_ups_1_d_payload_source,
  output wire [2:0]    io_ups_1_d_payload_size,
  output wire          io_ups_1_d_payload_denied,
  output wire [63:0]   io_ups_1_d_payload_data,
  output wire          io_ups_1_d_payload_corrupt,
  output wire          io_down_a_valid,
  input  wire          io_down_a_ready,
  output wire [2:0]    io_down_a_payload_opcode,
  output wire [2:0]    io_down_a_payload_param,
  output wire [1:0]    io_down_a_payload_source,
  output wire [31:0]   io_down_a_payload_address,
  output wire [2:0]    io_down_a_payload_size,
  output wire [7:0]    io_down_a_payload_mask,
  output wire [63:0]   io_down_a_payload_data,
  output wire          io_down_a_payload_corrupt,
  input  wire          io_down_d_valid,
  output wire          io_down_d_ready,
  input  wire [2:0]    io_down_d_payload_opcode,
  input  wire [2:0]    io_down_d_payload_param,
  input  wire [1:0]    io_down_d_payload_source,
  input  wire [2:0]    io_down_d_payload_size,
  input  wire          io_down_d_payload_denied,
  input  wire [63:0]   io_down_d_payload_data,
  input  wire          io_down_d_payload_corrupt,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire                a_arbiter_io_inputs_0_ready;
  wire                a_arbiter_io_inputs_1_ready;
  wire                a_arbiter_io_output_valid;
  wire       [2:0]    a_arbiter_io_output_payload_opcode;
  wire       [2:0]    a_arbiter_io_output_payload_param;
  wire       [1:0]    a_arbiter_io_output_payload_source;
  wire       [31:0]   a_arbiter_io_output_payload_address;
  wire       [2:0]    a_arbiter_io_output_payload_size;
  wire       [7:0]    a_arbiter_io_output_payload_mask;
  wire       [63:0]   a_arbiter_io_output_payload_data;
  wire                a_arbiter_io_output_payload_corrupt;
  wire       [0:0]    a_arbiter_io_chosen;
  wire       [1:0]    a_arbiter_io_chosenOH;
  wire       [1:0]    _zz_ups_1_a_payload_source;
  reg                 _zz_io_down_d_ready;
  wire                ups_0_a_valid;
  wire                ups_0_a_ready;
  wire       [2:0]    ups_0_a_payload_opcode;
  wire       [2:0]    ups_0_a_payload_param;
  wire       [1:0]    ups_0_a_payload_source;
  wire       [31:0]   ups_0_a_payload_address;
  wire       [2:0]    ups_0_a_payload_size;
  wire                ups_0_d_valid;
  wire                ups_0_d_ready;
  wire       [2:0]    ups_0_d_payload_opcode;
  wire       [2:0]    ups_0_d_payload_param;
  wire       [1:0]    ups_0_d_payload_source;
  wire       [2:0]    ups_0_d_payload_size;
  wire                ups_0_d_payload_denied;
  wire       [63:0]   ups_0_d_payload_data;
  wire                ups_0_d_payload_corrupt;
  wire                ups_1_a_valid;
  wire                ups_1_a_ready;
  wire       [2:0]    ups_1_a_payload_opcode;
  wire       [2:0]    ups_1_a_payload_param;
  wire       [1:0]    ups_1_a_payload_source;
  wire       [31:0]   ups_1_a_payload_address;
  wire       [2:0]    ups_1_a_payload_size;
  wire       [7:0]    ups_1_a_payload_mask;
  wire       [63:0]   ups_1_a_payload_data;
  wire                ups_1_a_payload_corrupt;
  wire                ups_1_d_valid;
  wire                ups_1_d_ready;
  wire       [2:0]    ups_1_d_payload_opcode;
  wire       [2:0]    ups_1_d_payload_param;
  wire       [1:0]    ups_1_d_payload_source;
  wire       [2:0]    ups_1_d_payload_size;
  wire                ups_1_d_payload_denied;
  wire       [63:0]   ups_1_d_payload_data;
  wire                ups_1_d_payload_corrupt;
  wire       [0:0]    d_sel;
  `ifndef SYNTHESIS
  reg [127:0] io_ups_0_a_payload_opcode_string;
  reg [119:0] io_ups_0_d_payload_opcode_string;
  reg [127:0] io_ups_1_a_payload_opcode_string;
  reg [119:0] io_ups_1_d_payload_opcode_string;
  reg [127:0] io_down_a_payload_opcode_string;
  reg [119:0] io_down_d_payload_opcode_string;
  reg [127:0] ups_0_a_payload_opcode_string;
  reg [119:0] ups_0_d_payload_opcode_string;
  reg [127:0] ups_1_a_payload_opcode_string;
  reg [119:0] ups_1_d_payload_opcode_string;
  `endif


  assign _zz_ups_1_a_payload_source = {1'd0, io_ups_1_a_payload_source};
  StreamArbiter_5 a_arbiter (
    .io_inputs_0_valid           (ups_0_a_valid                                                       ), //i
    .io_inputs_0_ready           (a_arbiter_io_inputs_0_ready                                         ), //o
    .io_inputs_0_payload_opcode  (ups_0_a_payload_opcode[2:0]                                         ), //i
    .io_inputs_0_payload_param   (ups_0_a_payload_param[2:0]                                          ), //i
    .io_inputs_0_payload_source  (ups_0_a_payload_source[1:0]                                         ), //i
    .io_inputs_0_payload_address (ups_0_a_payload_address[31:0]                                       ), //i
    .io_inputs_0_payload_size    (ups_0_a_payload_size[2:0]                                           ), //i
    .io_inputs_0_payload_mask    (8'bxxxxxxxx                                                         ), //i
    .io_inputs_0_payload_data    (64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx), //i
    .io_inputs_0_payload_corrupt (1'b0                                                                ), //i
    .io_inputs_1_valid           (ups_1_a_valid                                                       ), //i
    .io_inputs_1_ready           (a_arbiter_io_inputs_1_ready                                         ), //o
    .io_inputs_1_payload_opcode  (ups_1_a_payload_opcode[2:0]                                         ), //i
    .io_inputs_1_payload_param   (ups_1_a_payload_param[2:0]                                          ), //i
    .io_inputs_1_payload_source  (ups_1_a_payload_source[1:0]                                         ), //i
    .io_inputs_1_payload_address (ups_1_a_payload_address[31:0]                                       ), //i
    .io_inputs_1_payload_size    (ups_1_a_payload_size[2:0]                                           ), //i
    .io_inputs_1_payload_mask    (ups_1_a_payload_mask[7:0]                                           ), //i
    .io_inputs_1_payload_data    (ups_1_a_payload_data[63:0]                                          ), //i
    .io_inputs_1_payload_corrupt (ups_1_a_payload_corrupt                                             ), //i
    .io_output_valid             (a_arbiter_io_output_valid                                           ), //o
    .io_output_ready             (io_down_a_ready                                                     ), //i
    .io_output_payload_opcode    (a_arbiter_io_output_payload_opcode[2:0]                             ), //o
    .io_output_payload_param     (a_arbiter_io_output_payload_param[2:0]                              ), //o
    .io_output_payload_source    (a_arbiter_io_output_payload_source[1:0]                             ), //o
    .io_output_payload_address   (a_arbiter_io_output_payload_address[31:0]                           ), //o
    .io_output_payload_size      (a_arbiter_io_output_payload_size[2:0]                               ), //o
    .io_output_payload_mask      (a_arbiter_io_output_payload_mask[7:0]                               ), //o
    .io_output_payload_data      (a_arbiter_io_output_payload_data[63:0]                              ), //o
    .io_output_payload_corrupt   (a_arbiter_io_output_payload_corrupt                                 ), //o
    .io_chosen                   (a_arbiter_io_chosen                                                 ), //o
    .io_chosenOH                 (a_arbiter_io_chosenOH[1:0]                                          ), //o
    .litex_clk                   (litex_clk                                                           ), //i
    .cpuResetCtrl_reset          (cpuResetCtrl_reset                                                  )  //i
  );
  always @(*) begin
    case(d_sel)
      1'b0 : _zz_io_down_d_ready = ups_0_d_ready;
      default : _zz_io_down_d_ready = ups_1_d_ready;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_ups_0_a_payload_opcode)
      A_PUT_FULL_DATA : io_ups_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_ups_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_ups_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_ups_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_ups_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_ups_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_0_d_payload_opcode)
      D_ACCESS_ACK : io_ups_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_ups_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_ups_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_ups_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_ups_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_ups_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_1_a_payload_opcode)
      A_PUT_FULL_DATA : io_ups_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_ups_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_ups_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_ups_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_ups_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_ups_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_ups_1_d_payload_opcode)
      D_ACCESS_ACK : io_ups_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_ups_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_ups_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_ups_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_ups_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_ups_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_down_a_payload_opcode)
      A_PUT_FULL_DATA : io_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_down_d_payload_opcode)
      D_ACCESS_ACK : io_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : io_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ups_0_a_payload_opcode)
      A_PUT_FULL_DATA : ups_0_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ups_0_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ups_0_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ups_0_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ups_0_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ups_0_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ups_0_d_payload_opcode)
      D_ACCESS_ACK : ups_0_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ups_0_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ups_0_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ups_0_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ups_0_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ups_0_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(ups_1_a_payload_opcode)
      A_PUT_FULL_DATA : ups_1_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : ups_1_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : ups_1_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : ups_1_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : ups_1_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : ups_1_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(ups_1_d_payload_opcode)
      D_ACCESS_ACK : ups_1_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : ups_1_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : ups_1_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : ups_1_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : ups_1_d_payload_opcode_string = "RELEASE_ACK    ";
      default : ups_1_d_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign ups_0_a_valid = io_ups_0_a_valid;
  assign io_ups_0_a_ready = ups_0_a_ready;
  assign ups_0_a_payload_opcode = io_ups_0_a_payload_opcode;
  assign ups_0_a_payload_param = io_ups_0_a_payload_param;
  assign ups_0_a_payload_address = io_ups_0_a_payload_address;
  assign ups_0_a_payload_size = io_ups_0_a_payload_size;
  assign io_ups_0_d_valid = ups_0_d_valid;
  assign ups_0_d_ready = io_ups_0_d_ready;
  assign io_ups_0_d_payload_opcode = ups_0_d_payload_opcode;
  assign io_ups_0_d_payload_param = ups_0_d_payload_param;
  assign io_ups_0_d_payload_size = ups_0_d_payload_size;
  assign io_ups_0_d_payload_denied = ups_0_d_payload_denied;
  assign io_ups_0_d_payload_data = ups_0_d_payload_data;
  assign io_ups_0_d_payload_corrupt = ups_0_d_payload_corrupt;
  assign ups_0_a_payload_source = (2'b00 | 2'b00);
  assign ups_1_a_valid = io_ups_1_a_valid;
  assign io_ups_1_a_ready = ups_1_a_ready;
  assign ups_1_a_payload_opcode = io_ups_1_a_payload_opcode;
  assign ups_1_a_payload_param = io_ups_1_a_payload_param;
  assign ups_1_a_payload_address = io_ups_1_a_payload_address;
  assign ups_1_a_payload_size = io_ups_1_a_payload_size;
  assign ups_1_a_payload_mask = io_ups_1_a_payload_mask;
  assign ups_1_a_payload_data = io_ups_1_a_payload_data;
  assign ups_1_a_payload_corrupt = io_ups_1_a_payload_corrupt;
  assign io_ups_1_d_valid = ups_1_d_valid;
  assign ups_1_d_ready = io_ups_1_d_ready;
  assign io_ups_1_d_payload_opcode = ups_1_d_payload_opcode;
  assign io_ups_1_d_payload_param = ups_1_d_payload_param;
  assign io_ups_1_d_payload_size = ups_1_d_payload_size;
  assign io_ups_1_d_payload_denied = ups_1_d_payload_denied;
  assign io_ups_1_d_payload_data = ups_1_d_payload_data;
  assign io_ups_1_d_payload_corrupt = ups_1_d_payload_corrupt;
  assign ups_1_a_payload_source = (_zz_ups_1_a_payload_source | 2'b10);
  assign io_ups_1_d_payload_source = ups_1_d_payload_source[0:0];
  assign ups_0_a_ready = a_arbiter_io_inputs_0_ready;
  assign ups_1_a_ready = a_arbiter_io_inputs_1_ready;
  assign io_down_a_valid = a_arbiter_io_output_valid;
  assign io_down_a_payload_opcode = a_arbiter_io_output_payload_opcode;
  assign io_down_a_payload_param = a_arbiter_io_output_payload_param;
  assign io_down_a_payload_source = a_arbiter_io_output_payload_source;
  assign io_down_a_payload_address = a_arbiter_io_output_payload_address;
  assign io_down_a_payload_size = a_arbiter_io_output_payload_size;
  assign io_down_a_payload_mask = a_arbiter_io_output_payload_mask;
  assign io_down_a_payload_data = a_arbiter_io_output_payload_data;
  assign io_down_a_payload_corrupt = a_arbiter_io_output_payload_corrupt;
  assign d_sel = io_down_d_payload_source[1 : 1];
  assign io_down_d_ready = _zz_io_down_d_ready;
  assign ups_0_d_valid = (io_down_d_valid && (d_sel == 1'b0));
  assign ups_0_d_payload_opcode = io_down_d_payload_opcode;
  assign ups_0_d_payload_param = io_down_d_payload_param;
  assign ups_0_d_payload_source = io_down_d_payload_source;
  assign ups_0_d_payload_denied = io_down_d_payload_denied;
  assign ups_0_d_payload_size = io_down_d_payload_size;
  assign ups_0_d_payload_data = io_down_d_payload_data;
  assign ups_0_d_payload_corrupt = io_down_d_payload_corrupt;
  assign ups_1_d_valid = (io_down_d_valid && (d_sel == 1'b1));
  assign ups_1_d_payload_opcode = io_down_d_payload_opcode;
  assign ups_1_d_payload_param = io_down_d_payload_param;
  assign ups_1_d_payload_source = io_down_d_payload_source;
  assign ups_1_d_payload_denied = io_down_d_payload_denied;
  assign ups_1_d_payload_size = io_down_d_payload_size;
  assign ups_1_d_payload_data = io_down_d_payload_data;
  assign ups_1_d_payload_corrupt = io_down_d_payload_corrupt;

endmodule

module BufferCC_1 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_fiber_holder_reset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge litex_clk or posedge cpuResetCtrl_fiber_holder_reset) begin
    if(cpuResetCtrl_fiber_holder_reset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          litex_clk,
  input  wire          litex_reset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge litex_clk or posedge litex_reset) begin
    if(litex_reset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module VexiiRiscv (
  output wire          CfuPlugin_logic_bus_cmd_valid,
  input  wire          CfuPlugin_logic_bus_cmd_ready,
  output wire [2:0]    CfuPlugin_logic_bus_cmd_payload_function_id,
  output wire [31:0]   CfuPlugin_logic_bus_cmd_payload_inputs_0,
  output wire [31:0]   CfuPlugin_logic_bus_cmd_payload_inputs_1,
  output wire [2:0]    CfuPlugin_logic_bus_cmd_payload_state_index,
  output wire [3:0]    CfuPlugin_logic_bus_cmd_payload_cfu_index,
  output wire [31:0]   CfuPlugin_logic_bus_cmd_payload_raw_insn,
  input  wire          CfuPlugin_logic_bus_rsp_valid,
  output wire          CfuPlugin_logic_bus_rsp_ready,
  input  wire [31:0]   CfuPlugin_logic_bus_rsp_payload_outputs_0,
  input  wire [63:0]   PrivilegedPlugin_logic_rdtime,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_timer /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_software /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_m_external /* verilator public */ ,
  input  wire          PrivilegedPlugin_logic_harts_0_int_s_external /* verilator public */ ,
  output wire          FetchL1TileLinkPlugin_logic_down_a_valid,
  input  wire          FetchL1TileLinkPlugin_logic_down_a_ready,
  output wire [2:0]    FetchL1TileLinkPlugin_logic_down_a_payload_opcode,
  output wire [2:0]    FetchL1TileLinkPlugin_logic_down_a_payload_param,
  output wire [31:0]   FetchL1TileLinkPlugin_logic_down_a_payload_address,
  output wire [2:0]    FetchL1TileLinkPlugin_logic_down_a_payload_size,
  input  wire          FetchL1TileLinkPlugin_logic_down_d_valid,
  output wire          FetchL1TileLinkPlugin_logic_down_d_ready,
  input  wire [2:0]    FetchL1TileLinkPlugin_logic_down_d_payload_opcode,
  input  wire [2:0]    FetchL1TileLinkPlugin_logic_down_d_payload_param,
  input  wire [2:0]    FetchL1TileLinkPlugin_logic_down_d_payload_size,
  input  wire          FetchL1TileLinkPlugin_logic_down_d_payload_denied,
  input  wire [63:0]   FetchL1TileLinkPlugin_logic_down_d_payload_data,
  input  wire          FetchL1TileLinkPlugin_logic_down_d_payload_corrupt,
  output reg           LsuL1TileLinkPlugin_logic_down_a_valid,
  input  wire          LsuL1TileLinkPlugin_logic_down_a_ready,
  output reg  [2:0]    LsuL1TileLinkPlugin_logic_down_a_payload_opcode,
  output wire [2:0]    LsuL1TileLinkPlugin_logic_down_a_payload_param,
  output reg  [0:0]    LsuL1TileLinkPlugin_logic_down_a_payload_source,
  output reg  [31:0]   LsuL1TileLinkPlugin_logic_down_a_payload_address,
  output wire [2:0]    LsuL1TileLinkPlugin_logic_down_a_payload_size,
  output wire [7:0]    LsuL1TileLinkPlugin_logic_down_a_payload_mask,
  output wire [63:0]   LsuL1TileLinkPlugin_logic_down_a_payload_data,
  output wire          LsuL1TileLinkPlugin_logic_down_a_payload_corrupt,
  input  wire          LsuL1TileLinkPlugin_logic_down_d_valid,
  output wire          LsuL1TileLinkPlugin_logic_down_d_ready,
  input  wire [2:0]    LsuL1TileLinkPlugin_logic_down_d_payload_opcode,
  input  wire [2:0]    LsuL1TileLinkPlugin_logic_down_d_payload_param,
  input  wire [0:0]    LsuL1TileLinkPlugin_logic_down_d_payload_source,
  input  wire [2:0]    LsuL1TileLinkPlugin_logic_down_d_payload_size,
  input  wire          LsuL1TileLinkPlugin_logic_down_d_payload_denied,
  input  wire [63:0]   LsuL1TileLinkPlugin_logic_down_d_payload_data,
  input  wire          LsuL1TileLinkPlugin_logic_down_d_payload_corrupt,
  output wire          LsuTileLinkPlugin_logic_bridge_down_a_valid,
  input  wire          LsuTileLinkPlugin_logic_bridge_down_a_ready,
  output wire [2:0]    LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode,
  output wire [2:0]    LsuTileLinkPlugin_logic_bridge_down_a_payload_param,
  output wire [31:0]   LsuTileLinkPlugin_logic_bridge_down_a_payload_address,
  output wire [1:0]    LsuTileLinkPlugin_logic_bridge_down_a_payload_size,
  output wire [3:0]    LsuTileLinkPlugin_logic_bridge_down_a_payload_mask,
  output wire [31:0]   LsuTileLinkPlugin_logic_bridge_down_a_payload_data,
  output wire          LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt,
  input  wire          LsuTileLinkPlugin_logic_bridge_down_d_valid,
  output wire          LsuTileLinkPlugin_logic_bridge_down_d_ready,
  input  wire [2:0]    LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode,
  input  wire [2:0]    LsuTileLinkPlugin_logic_bridge_down_d_payload_param,
  input  wire [1:0]    LsuTileLinkPlugin_logic_bridge_down_d_payload_size,
  input  wire          LsuTileLinkPlugin_logic_bridge_down_d_payload_denied,
  input  wire [31:0]   LsuTileLinkPlugin_logic_bridge_down_d_payload_data,
  input  wire          LsuTileLinkPlugin_logic_bridge_down_d_payload_corrupt,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);
  localparam BranchPlugin_BranchCtrlEnum_B = 2'd0;
  localparam BranchPlugin_BranchCtrlEnum_JAL = 2'd1;
  localparam BranchPlugin_BranchCtrlEnum_JALR = 2'd2;
  localparam EnvPluginOp_ECALL = 3'd0;
  localparam EnvPluginOp_EBREAK = 3'd1;
  localparam EnvPluginOp_PRIV_RET = 3'd2;
  localparam EnvPluginOp_FENCE_I = 3'd3;
  localparam EnvPluginOp_SFENCE_VMA = 3'd4;
  localparam EnvPluginOp_WFI = 3'd5;
  localparam Input2Kind_RS = 1'd0;
  localparam Input2Kind_IMM_I = 1'd1;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 = 2'd0;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_OR_1 = 2'd1;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_AND_1 = 2'd2;
  localparam IntAluPlugin_AluBitwiseCtrlEnum_ZERO = 2'd3;
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;
  localparam TrapPlugin_logic_harts_0_trap_fsm_RESET = 4'd0;
  localparam TrapPlugin_logic_harts_0_trap_fsm_RUNNING = 4'd1;
  localparam TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 = 4'd2;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC = 4'd3;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL = 4'd4;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC = 4'd5;
  localparam TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY = 4'd6;
  localparam TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC = 4'd7;
  localparam TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY = 4'd8;
  localparam TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP = 4'd9;
  localparam TrapPlugin_logic_harts_0_trap_fsm_JUMP = 4'd10;
  localparam TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH = 4'd11;
  localparam TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH = 4'd12;
  localparam LsuL1CmdOpcode_LSU = 3'd0;
  localparam LsuL1CmdOpcode_ACCESS_1 = 3'd1;
  localparam LsuL1CmdOpcode_STORE_BUFFER = 3'd2;
  localparam LsuL1CmdOpcode_FLUSH = 3'd3;
  localparam LsuL1CmdOpcode_PREFETCH = 3'd4;
  localparam LsuPlugin_logic_flusher_IDLE = 2'd0;
  localparam LsuPlugin_logic_flusher_CMD = 2'd1;
  localparam LsuPlugin_logic_flusher_COMPLETION = 2'd2;
  localparam MmuPlugin_logic_refill_BOOT = 3'd0;
  localparam MmuPlugin_logic_refill_IDLE = 3'd1;
  localparam MmuPlugin_logic_refill_CMD_0 = 3'd2;
  localparam MmuPlugin_logic_refill_CMD_1 = 3'd3;
  localparam MmuPlugin_logic_refill_RSP_0 = 3'd4;
  localparam MmuPlugin_logic_refill_RSP_1 = 3'd5;
  localparam CsrAccessPlugin_logic_fsm_IDLE = 2'd0;
  localparam CsrAccessPlugin_logic_fsm_READ = 2'd1;
  localparam CsrAccessPlugin_logic_fsm_WRITE = 2'd2;
  localparam CsrAccessPlugin_logic_fsm_COMPLETION = 2'd3;
  localparam PerformanceCounterPlugin_logic_fsm_BOOT = 3'd0;
  localparam PerformanceCounterPlugin_logic_fsm_IDLE = 3'd1;
  localparam PerformanceCounterPlugin_logic_fsm_READ_LOW = 3'd2;
  localparam PerformanceCounterPlugin_logic_fsm_CALC_LOW = 3'd3;
  localparam PerformanceCounterPlugin_logic_fsm_READ_HIGH = 3'd4;
  localparam PerformanceCounterPlugin_logic_fsm_CALC_HIGH = 3'd5;
  localparam PerformanceCounterPlugin_logic_fsm_CSR_WRITE = 3'd6;

  wire                early0_DivPlugin_logic_processing_div_io_cmd_valid;
  wire                CfuPlugin_logic_onJoin_busRspStream_fifo_io_pop_ready;
  reg                 LsuPlugin_logic_flusher_arbiter_io_output_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_ready;
  reg                 MmuPlugin_logic_refill_arbiter_io_output_ready;
  reg                 MmuPlugin_logic_invalidate_arbiter_io_output_ready;
  reg                 integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid;
  reg        [4:0]    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address;
  reg        [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data;
  wire                BtbPlugin_logic_ras_mem_stack_wr_en;
  wire       [29:0]   BtbPlugin_logic_ras_mem_stack_wr_data;
  wire                LsuL1Plugin_logic_banks_0_mem_wr_en;
  wire                LsuL1Plugin_logic_banks_0_mem_rd_en;
  wire                LsuL1Plugin_logic_banks_1_mem_wr_en;
  wire                LsuL1Plugin_logic_banks_1_mem_rd_en;
  wire                LsuL1Plugin_logic_banks_2_mem_wr_en;
  wire                LsuL1Plugin_logic_banks_2_mem_rd_en;
  wire                LsuL1Plugin_logic_banks_3_mem_wr_en;
  wire                LsuL1Plugin_logic_banks_3_mem_rd_en;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_wr_en;
  wire       [39:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_wr_data;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_wr_en;
  wire       [39:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_wr_data;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_wr_en;
  wire       [19:0]   FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_wr_data;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_wr_en;
  wire       [39:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_wr_data;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_wr_en;
  wire       [39:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_wr_data;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_wr_en;
  wire       [39:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_wr_data;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_wr_en;
  wire       [19:0]   LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_wr_data;
  reg        [63:0]   FetchL1Plugin_logic_banks_0_mem_spinal_port1;
  reg        [63:0]   FetchL1Plugin_logic_banks_1_mem_spinal_port1;
  reg        [63:0]   FetchL1Plugin_logic_banks_2_mem_spinal_port1;
  reg        [63:0]   FetchL1Plugin_logic_banks_3_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_0_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_1_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_2_mem_spinal_port1;
  reg        [21:0]   FetchL1Plugin_logic_ways_3_mem_spinal_port1;
  reg        [2:0]    FetchL1Plugin_logic_plru_mem_spinal_port1;
  reg        [1:0]    GSharePlugin_logic_mem_counter_spinal_port1;
  reg        [48:0]   BtbPlugin_logic_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_0_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_1_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_2_mem_spinal_port1;
  reg        [21:0]   LsuL1Plugin_logic_ways_3_mem_spinal_port1;
  reg        [6:0]    LsuL1Plugin_logic_shared_mem_spinal_port1;
  reg        [63:0]   LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1;
  reg        [31:0]   CsrRamPlugin_logic_mem_spinal_port1;
  wire                early0_DivPlugin_logic_processing_div_io_cmd_ready;
  wire                early0_DivPlugin_logic_processing_div_io_rsp_valid;
  wire       [31:0]   early0_DivPlugin_logic_processing_div_io_rsp_payload_result;
  wire       [31:0]   early0_DivPlugin_logic_processing_div_io_rsp_payload_remain;
  wire                CfuPlugin_logic_onJoin_busRspStream_fifo_io_push_ready;
  wire                CfuPlugin_logic_onJoin_busRspStream_fifo_io_pop_valid;
  wire       [31:0]   CfuPlugin_logic_onJoin_busRspStream_fifo_io_pop_payload_outputs_0;
  wire       [1:0]    CfuPlugin_logic_onJoin_busRspStream_fifo_io_occupancy;
  wire       [1:0]    CfuPlugin_logic_onJoin_busRspStream_fifo_io_availability;
  wire                LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready;
  wire                LsuPlugin_logic_flusher_arbiter_io_output_valid;
  wire       [0:0]    LsuPlugin_logic_flusher_arbiter_io_chosenOH;
  wire                streamArbiter_10_io_inputs_0_ready;
  wire                streamArbiter_10_io_output_valid;
  wire       [31:0]   streamArbiter_10_io_output_payload_pcOnLastSlice;
  wire       [31:0]   streamArbiter_10_io_output_payload_pcTarget;
  wire                streamArbiter_10_io_output_payload_taken;
  wire                streamArbiter_10_io_output_payload_isBranch;
  wire                streamArbiter_10_io_output_payload_isPush;
  wire                streamArbiter_10_io_output_payload_isPop;
  wire                streamArbiter_10_io_output_payload_wasWrong;
  wire                streamArbiter_10_io_output_payload_badPredictedTarget;
  wire       [11:0]   streamArbiter_10_io_output_payload_history;
  wire       [15:0]   streamArbiter_10_io_output_payload_uopId;
  wire       [1:0]    streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire       [0:0]    streamArbiter_10_io_chosenOH;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_valid;
  wire       [2:0]    LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_clean;
  wire                LsuPlugin_logic_onAddress0_arbiter_io_output_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId;
  wire       [1:0]    LsuPlugin_logic_onAddress0_arbiter_io_chosen;
  wire       [2:0]    LsuPlugin_logic_onAddress0_arbiter_io_chosenOH;
  wire                MmuPlugin_logic_refill_arbiter_io_inputs_0_ready;
  wire                MmuPlugin_logic_refill_arbiter_io_output_valid;
  wire       [31:0]   MmuPlugin_logic_refill_arbiter_io_output_payload_address;
  wire       [0:0]    MmuPlugin_logic_refill_arbiter_io_output_payload_storageId;
  wire       [0:0]    MmuPlugin_logic_refill_arbiter_io_chosenOH;
  wire                MmuPlugin_logic_invalidate_arbiter_io_inputs_0_ready;
  wire                MmuPlugin_logic_invalidate_arbiter_io_output_valid;
  wire       [0:0]    MmuPlugin_logic_invalidate_arbiter_io_chosenOH;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  wire       [31:0]   integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  wire       [29:0]   BtbPlugin_logic_ras_mem_stack_rd_data;
  wire       [63:0]   LsuL1Plugin_logic_banks_0_mem_rd_data;
  wire       [63:0]   LsuL1Plugin_logic_banks_1_mem_rd_data;
  wire       [63:0]   LsuL1Plugin_logic_banks_2_mem_rd_data;
  wire       [63:0]   LsuL1Plugin_logic_banks_3_mem_rd_data;
  wire       [39:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_rd_data;
  wire       [39:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_rd_data;
  wire       [19:0]   FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_rd_data;
  wire       [39:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_rd_data;
  wire       [39:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_rd_data;
  wire       [39:0]   LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_rd_data;
  wire       [19:0]   LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_rd_data;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_1;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_2;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_3;
  wire       [31:0]   _zz_early0_IntAluPlugin_logic_alu_result_4;
  wire       [0:0]    _zz_early0_IntAluPlugin_logic_alu_result_5;
  wire       [4:0]    _zz_early0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_1;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_2;
  wire       [20:0]   _zz_early0_BarrelShifterPlugin_logic_shift_reversed_3;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_reversed_4;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_5;
  wire       [9:0]    _zz_early0_BarrelShifterPlugin_logic_shift_reversed_6;
  wire       [32:0]   _zz_early0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [32:0]   _zz_early0_BarrelShifterPlugin_logic_shift_shifted_1;
  wire       [31:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_1;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_2;
  wire       [20:0]   _zz_early0_BarrelShifterPlugin_logic_shift_patched_3;
  wire                _zz_early0_BarrelShifterPlugin_logic_shift_patched_4;
  wire       [0:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_5;
  wire       [9:0]    _zz_early0_BarrelShifterPlugin_logic_shift_patched_6;
  wire       [32:0]   _zz_execute_ctrl2_down_MUL_SRC1_lane0;
  wire       [32:0]   _zz_execute_ctrl2_down_MUL_SRC2_lane0;
  wire       [46:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_1;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_2;
  wire       [15:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_3;
  wire       [46:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [33:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_1;
  wire       [15:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_2;
  wire       [17:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_3;
  wire       [29:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_1;
  wire       [15:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_2;
  wire       [15:0]   _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_3;
  wire       [62:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3;
  wire       [62:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4;
  wire       [62:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5;
  wire       [62:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6;
  wire       [4:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3;
  wire       [4:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4;
  wire       [4:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5;
  wire       [4:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6;
  wire       [31:0]   _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2;
  wire       [0:0]    _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_0_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_0_mem_port_1;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_1_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_1_mem_port_1;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_2_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_2_mem_port_1;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_3_mem_port;
  wire                _zz_FetchL1Plugin_logic_ways_3_mem_port_1;
  wire       [2:0]    _zz_FetchL1Plugin_logic_plru_mem_port;
  wire                _zz_when;
  reg        [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [0:0]    _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0_1;
  reg        [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire       [0:0]    _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1_1;
  reg        [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2;
  wire       [0:0]    _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2_1;
  reg        [31:0]   _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3;
  wire       [0:0]    _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3_1;
  wire       [19:0]   _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits;
  wire       [19:0]   _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits;
  wire       [19:0]   _zz_FetchL1Plugin_logic_hits_w_2_indirect_bypassHits;
  wire       [19:0]   _zz_FetchL1Plugin_logic_hits_w_3_indirect_bypassHits;
  wire       [0:0]    _zz_FetchL1Plugin_logic_ctrl_dataAccessFault;
  wire       [1:0]    _zz_GSharePlugin_logic_mem_counter_port;
  wire                _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1;
  wire       [0:0]    _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2;
  wire       [5:0]    _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_3;
  wire       [13:0]   _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_4;
  wire       [11:0]   _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_5;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push_1;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_push_2;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_push_3;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_push_4;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2;
  wire       [1:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3;
  wire       [0:0]    _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4;
  wire       [48:0]   _zz_BtbPlugin_logic_mem_port;
  wire       [63:0]   _zz_WhiteboxerPlugin_logic_decodes_0_pc;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_commitCount;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_commitCount_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_eventInstructions_0;
  wire       [7:0]    _zz_PerformanceCounterPlugin_logic_counters_cycle_value;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_counters_cycle_value_1;
  wire       [7:0]    _zz_PerformanceCounterPlugin_logic_counters_instret_value_1;
  wire       [11:0]   _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  wire       [11:0]   _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3;
  wire       [20:0]   _zz_early0_BranchPlugin_pcCalc_target_b;
  wire       [11:0]   _zz_early0_BranchPlugin_pcCalc_target_b_1;
  wire       [12:0]   _zz_early0_BranchPlugin_pcCalc_target_b_2;
  wire       [1:0]    _zz_early0_BranchPlugin_pcCalc_slices;
  wire       [0:0]    _zz_early0_BranchPlugin_pcCalc_slices_1;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  wire       [3:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1;
  wire       [31:0]   _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  wire       [1:0]    _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1;
  reg        [2:0]    _zz_CfuPlugin_logic_bus_cmd_payload_function_id;
  wire       [31:0]   _zz__zz_CfuPlugin_logic_bus_cmd_payload_inputs_1;
  wire       [7:0]    _zz__zz_CfuPlugin_logic_bus_cmd_payload_inputs_1_1;
  wire       [3:0]    _zz_early0_EnvPlugin_logic_trapPort_payload_code;
  wire       [31:0]   _zz_early0_BranchPlugin_logic_alu_expectedMsb;
  wire       [12:0]   _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS1_ENABLE_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_RS2_ENABLE_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS2_ENABLE_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RS2_ENABLE_0_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_2;
  wire       [31:0]   _zz_decode_ctrls_1_down_RD_ENABLE_0_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_0_4;
  wire       [0:0]    _zz_decode_ctrls_1_down_RD_ENABLE_0_5;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_1;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_2;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_4;
  wire       [18:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_5;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_6;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_7;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_8;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_9;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_10;
  wire       [12:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_11;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_12;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_13;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_14;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_15;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_16;
  wire       [6:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_17;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_18;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_19;
  wire       [31:0]   _zz_decode_ctrls_1_down_Decode_LEGAL_0_20;
  wire                _zz_decode_ctrls_1_down_Decode_LEGAL_0_21;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_22;
  wire       [0:0]    _zz_decode_ctrls_1_down_Decode_LEGAL_0_23;
  wire       [0:0]    _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb;
  wire       [31:0]   _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice;
  wire       [1:0]    _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress_1;
  wire                _zz_CsrRamPlugin_csrMapper_ramAddress_2;
  wire                _zz_CsrRamPlugin_csrMapper_ramAddress_3;
  wire                _zz_CsrRamPlugin_csrMapper_ramAddress_4;
  wire                _zz_CsrRamPlugin_csrMapper_ramAddress_5;
  wire                _zz_GSharePlugin_logic_onLearn_hash_1;
  wire       [0:0]    _zz_GSharePlugin_logic_onLearn_hash_2;
  wire       [5:0]    _zz_GSharePlugin_logic_onLearn_hash_3;
  wire       [13:0]   _zz_GSharePlugin_logic_onLearn_hash_4;
  wire       [11:0]   _zz_GSharePlugin_logic_onLearn_hash_5;
  wire       [29:0]   _zz_BtbPlugin_logic_memWrite_payload_address;
  wire       [0:0]    _zz_decode_ctrls_1_down_CfuPlugin_logic_CFU_ENABLE_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_CfuPlugin_logic_CFU_ENABLE_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_2;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3;
  wire       [0:0]    _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_4;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1;
  wire       [0:0]    _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_2;
  wire       [29:0]   _zz_BtbPlugin_logic_memWrite_payload_address_1;
  wire       [29:0]   _zz_BtbPlugin_logic_memRead_cmd_payload;
  wire       [31:0]   _zz_BtbPlugin_logic_ras_write_payload_data;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_0_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_0_mem_port_1;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_1_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_1_mem_port_1;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_2_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_2_mem_port_1;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_3_mem_port;
  wire                _zz_LsuL1Plugin_logic_ways_3_mem_port_1;
  wire       [6:0]    _zz_LsuL1Plugin_logic_shared_mem_port;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_read_wordIndex;
  wire       [0:0]    _zz_LsuL1Plugin_logic_writeback_read_wordIndex_1;
  reg        [63:0]   _zz_LsuL1Plugin_logic_writeback_read_readedData;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_victimBuffer_port;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_write_wordIndex;
  wire       [0:0]    _zz_LsuL1Plugin_logic_writeback_write_wordIndex_1;
  reg        [31:0]   _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [0:0]    _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0_1;
  reg        [31:0]   _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [0:0]    _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1_1;
  reg        [31:0]   _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2;
  wire       [0:0]    _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2_1;
  reg        [31:0]   _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3;
  wire       [0:0]    _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3_1;
  wire       [3:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback;
  wire       [0:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_doWrite;
  wire       [2:0]    _zz_58;
  reg        [2:0]    _zz_59;
  wire       [2:0]    _zz_60;
  reg        [2:0]    _zz_61;
  wire       [2:0]    _zz_62;
  wire       [0:0]    _zz_63;
  reg        [1:0]    _zz_64;
  wire       [2:0]    _zz_65;
  wire       [3:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty_1;
  reg        [19:0]   _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address;
  reg                 _zz_LsuL1Plugin_logic_waysWrite_tag_fault;
  reg        [19:0]   _zz_LsuL1Plugin_logic_writeback_push_payload_address;
  wire       [36:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  wire       [36:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1;
  wire       [36:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2;
  wire       [36:0]   _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3;
  wire       [0:0]    _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_4;
  wire       [31:0]   _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
  wire       [2:0]    _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_ls_storeId;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_ls_storeId_1;
  wire       [12:0]   _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_addressExtension;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted;
  wire       [1:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_1;
  reg        [7:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2;
  wire       [0:0]    _zz_LsuPlugin_logic_onCtrl_loadData_shifted_3;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3;
  wire       [31:0]   _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4;
  wire       [1:0]    _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5;
  wire       [5:0]    _zz_LsuPlugin_logic_onCtrl_rva_lrsc_age;
  wire       [0:0]    _zz_LsuPlugin_logic_onCtrl_rva_lrsc_age_1;
  wire       [2:0]    _zz_LsuPlugin_logic_trapPort_payload_code;
  wire       [5:0]    _zz_LsuPlugin_logic_flusher_cmdCounter;
  reg        [2:0]    _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last;
  wire       [31:0]   _zz_PcPlugin_logic_harts_0_self_pc;
  wire       [2:0]    _zz_PcPlugin_logic_harts_0_self_pc_1;
  wire       [0:0]    _zz_PcPlugin_logic_harts_0_aggregator_fault;
  wire       [0:0]    _zz_PcPlugin_logic_harts_0_aggregator_fault_1_1;
  wire       [1:0]    _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
  wire       [0:0]    _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext_1;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_4;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser;
  wire       [19:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_1;
  wire       [19:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_2;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_3;
  wire       [19:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_4;
  wire       [11:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_5;
  wire       [9:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_6;
  wire       [21:0]   _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_7;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_3;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire       [0:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire       [11:0]   _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated;
  wire       [11:0]   _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated_1;
  wire                _zz_fetch_logic_flushes_0_doIt;
  wire                _zz_fetch_logic_flushes_0_doIt_1;
  wire                _zz_fetch_logic_flushes_0_doIt_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_0_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_0_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_1_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_1_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_2_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_2_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_3_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_3_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_4_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_4_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_5_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_5_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_6_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_6_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_7_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_7_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_8_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_8_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_9_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_9_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_10_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_10_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_11_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_11_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_12_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_12_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_13_1;
  wire       [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_13_2;
  wire       [6:0]    _zz_PerformanceCounterPlugin_logic_fsm_calc_a;
  wire       [7:0]    _zz_PerformanceCounterPlugin_logic_fsm_calc_b;
  wire       [32:0]   _zz_PerformanceCounterPlugin_logic_fsm_calc_sum;
  wire       [8:0]    _zz_PerformanceCounterPlugin_logic_fsm_calc_sum_1;
  wire       [1:0]    _zz_PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked;
  wire       [11:0]   _zz_COMB_CSR_;
  wire                _zz_COMB_CSR__1;
  wire       [0:0]    _zz_COMB_CSR__2;
  wire       [166:0]  _zz_COMB_CSR__3;
  wire       [11:0]   _zz_COMB_CSR__4;
  wire                _zz_COMB_CSR__5;
  wire       [0:0]    _zz_COMB_CSR__6;
  wire       [158:0]  _zz_COMB_CSR__7;
  wire       [11:0]   _zz_COMB_CSR__8;
  wire                _zz_COMB_CSR__9;
  wire       [0:0]    _zz_COMB_CSR__10;
  wire       [150:0]  _zz_COMB_CSR__11;
  wire       [11:0]   _zz_COMB_CSR__12;
  wire                _zz_COMB_CSR__13;
  wire       [0:0]    _zz_COMB_CSR__14;
  wire       [142:0]  _zz_COMB_CSR__15;
  wire       [11:0]   _zz_COMB_CSR__16;
  wire                _zz_COMB_CSR__17;
  wire       [0:0]    _zz_COMB_CSR__18;
  wire       [134:0]  _zz_COMB_CSR__19;
  wire       [11:0]   _zz_COMB_CSR__20;
  wire                _zz_COMB_CSR__21;
  wire       [0:0]    _zz_COMB_CSR__22;
  wire       [126:0]  _zz_COMB_CSR__23;
  wire       [11:0]   _zz_COMB_CSR__24;
  wire                _zz_COMB_CSR__25;
  wire       [0:0]    _zz_COMB_CSR__26;
  wire       [118:0]  _zz_COMB_CSR__27;
  wire       [11:0]   _zz_COMB_CSR__28;
  wire                _zz_COMB_CSR__29;
  wire       [0:0]    _zz_COMB_CSR__30;
  wire       [110:0]  _zz_COMB_CSR__31;
  wire       [11:0]   _zz_COMB_CSR__32;
  wire                _zz_COMB_CSR__33;
  wire       [0:0]    _zz_COMB_CSR__34;
  wire       [102:0]  _zz_COMB_CSR__35;
  wire       [11:0]   _zz_COMB_CSR__36;
  wire                _zz_COMB_CSR__37;
  wire       [0:0]    _zz_COMB_CSR__38;
  wire       [94:0]   _zz_COMB_CSR__39;
  wire       [11:0]   _zz_COMB_CSR__40;
  wire                _zz_COMB_CSR__41;
  wire       [0:0]    _zz_COMB_CSR__42;
  wire       [86:0]   _zz_COMB_CSR__43;
  wire       [11:0]   _zz_COMB_CSR__44;
  wire                _zz_COMB_CSR__45;
  wire       [0:0]    _zz_COMB_CSR__46;
  wire       [78:0]   _zz_COMB_CSR__47;
  wire       [11:0]   _zz_COMB_CSR__48;
  wire                _zz_COMB_CSR__49;
  wire       [0:0]    _zz_COMB_CSR__50;
  wire       [70:0]   _zz_COMB_CSR__51;
  wire       [11:0]   _zz_COMB_CSR__52;
  wire                _zz_COMB_CSR__53;
  wire       [0:0]    _zz_COMB_CSR__54;
  wire       [62:0]   _zz_COMB_CSR__55;
  wire       [11:0]   _zz_COMB_CSR__56;
  wire                _zz_COMB_CSR__57;
  wire       [0:0]    _zz_COMB_CSR__58;
  wire       [54:0]   _zz_COMB_CSR__59;
  wire       [11:0]   _zz_COMB_CSR__60;
  wire                _zz_COMB_CSR__61;
  wire       [0:0]    _zz_COMB_CSR__62;
  wire       [46:0]   _zz_COMB_CSR__63;
  wire       [11:0]   _zz_COMB_CSR__64;
  wire                _zz_COMB_CSR__65;
  wire       [0:0]    _zz_COMB_CSR__66;
  wire       [38:0]   _zz_COMB_CSR__67;
  wire       [11:0]   _zz_COMB_CSR__68;
  wire                _zz_COMB_CSR__69;
  wire       [0:0]    _zz_COMB_CSR__70;
  wire       [30:0]   _zz_COMB_CSR__71;
  wire       [11:0]   _zz_COMB_CSR__72;
  wire                _zz_COMB_CSR__73;
  wire       [0:0]    _zz_COMB_CSR__74;
  wire       [22:0]   _zz_COMB_CSR__75;
  wire       [11:0]   _zz_COMB_CSR__76;
  wire                _zz_COMB_CSR__77;
  wire       [0:0]    _zz_COMB_CSR__78;
  wire       [14:0]   _zz_COMB_CSR__79;
  wire       [11:0]   _zz_COMB_CSR__80;
  wire                _zz_COMB_CSR__81;
  wire       [0:0]    _zz_COMB_CSR__82;
  wire       [6:0]    _zz_COMB_CSR__83;
  wire       [11:0]   _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
  wire                _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_1;
  wire       [0:0]    _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_2;
  wire       [6:0]    _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_3;
  wire       [11:0]   _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter;
  wire       [11:0]   _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_1;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_inject_implemented_1;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented_2;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_inject_implemented_3;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24;
  wire       [18:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29;
  wire       [18:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34;
  wire       [19:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38;
  wire       [18:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56;
  wire       [12:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_57;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_58;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_59;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_60;
  wire       [17:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_61;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_62;
  wire       [14:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_63;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_64;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_65;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_66;
  wire       [22:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_67;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_68;
  wire       [20:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_69;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_70;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_71;
  wire       [21:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_72;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_73;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_74;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_75;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_76;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_77;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_78;
  wire       [11:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_79;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_80;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_81;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_82;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_83;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_84;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_85;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_86;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_87;
  wire       [11:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_88;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_89;
  wire       [7:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_90;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_91;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_92;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_93;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_94;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_95;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_96;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_97;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_98;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_99;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_100;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_101;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_102;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_103;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_104;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_105;
  wire       [12:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_106;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_107;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_108;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_109;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_110;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_111;
  wire       [15:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_112;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_113;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_114;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_115;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_116;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_117;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_118;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_119;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_120;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_121;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_122;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_123;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_124;
  wire       [3:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_125;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_126;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_127;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_128;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_129;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_130;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_131;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_132;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_133;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_134;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_135;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_136;
  wire       [8:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_137;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_138;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_139;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_140;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_141;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_142;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_143;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_144;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_145;
  wire       [14:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_146;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_147;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_148;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_149;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_150;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_151;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_152;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_153;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_154;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_155;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_156;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_157;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_158;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_159;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_160;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_161;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_162;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_163;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_164;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_165;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_166;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_167;
  wire       [9:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_168;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_169;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_170;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_171;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_172;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_173;
  wire       [5:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_174;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_175;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_176;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_177;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_178;
  wire       [1:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_179;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_180;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_181;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_182;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_183;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_184;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_185;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_186;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_187;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_188;
  wire       [0:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_189;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_190;
  wire       [2:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_191;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_192;
  wire       [2:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_193;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_194;
  wire       [2:0]    _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_195;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_196;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_197;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_198;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_199;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_200;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_201;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_202;
  wire       [13:0]   _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_203;
  wire       [31:0]   _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [4:0]    _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1;
  wire       [0:0]    _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit;
  wire       [31:0]   _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault;
  wire       [31:0]   _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault_1;
  wire       [0:0]    _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io_1;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_cached_rsp_fault;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_cached_rsp_fault_1;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_cached_rsp_fault_2;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_cached_rsp_fault_3;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_cached_rsp_fault_4;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_cached_rsp_io_1;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit;
  wire       [0:0]    _zz_LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_io_rsp_fault;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_io_rsp_fault_1;
  wire       [31:0]   _zz_LsuPlugin_logic_onPma_io_rsp_fault_2;
  wire                _zz_LsuPlugin_logic_onPma_io_rsp_fault_3;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_io_rsp_fault_4;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_io_rsp_fault_5;
  wire       [0:0]    _zz_LsuPlugin_logic_onPma_io_rsp_io_1;
  wire       [3:0]    _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [2:0]    _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  reg        [3:0]    _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload;
  wire       [4:0]    _zz_CsrRamPlugin_logic_flush_counter;
  wire       [0:0]    _zz_CsrRamPlugin_logic_flush_counter_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_2;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_3;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_5;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_6;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_1;
  wire       [31:0]   _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_3;
  wire       [0:0]    _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_4;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_DivPlugin_REM_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_DivPlugin_REM_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_1;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_2;
  wire       [31:0]   _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_3;
  wire                _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_4;
  wire                _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_5;
  wire                _zz_when_ExecuteLanePlugin_l306_2;
  wire       [31:0]   _zz_WhiteboxerPlugin_logic_csr_access_payload_address;
  reg        [0:0]    _zz_WhiteboxerPlugin_logic_perf_candidatesCount;
  wire       [0:0]    _zz_WhiteboxerPlugin_logic_perf_candidatesCount_1;
  reg        [0:0]    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  wire       [0:0]    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1;
  wire       [59:0]   _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
  wire       [0:0]    _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1;
  wire       [1:0]    _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask;
  wire       [3:0]    _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask;
  wire       [3:0]    _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask_1;
  wire       [32:0]   _zz_PerformanceCounterPlugin_logic_writePort_data;
  wire       [32:0]   _zz_PerformanceCounterPlugin_logic_writePort_data_1;
  wire       [31:0]   _zz_PerformanceCounterPlugin_logic_counters_cycle_value_2;
  wire       [31:0]   _zz_PerformanceCounterPlugin_logic_counters_instret_value_2;
  wire                fetch_logic_ctrls_0_up_isReady;
  wire                fetch_logic_ctrls_0_up_isValid;
  reg        [31:0]   execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  reg                 execute_ctrl5_up_COMMIT_lane0;
  reg        [4:0]    execute_ctrl5_up_RD_PHYS_lane0;
  wire       [11:0]   execute_ctrl3_down_Decode_STORE_ID_lane0;
  wire                execute_ctrl3_down_LsuL1_PREFETCH_lane0;
  wire                execute_ctrl3_down_LsuL1_INVALID_lane0;
  wire                execute_ctrl3_down_LsuL1_CLEAN_lane0;
  wire       [3:0]    execute_ctrl3_down_LsuL1_MASK_lane0;
  wire                execute_ctrl3_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl3_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl3_down_AguPlugin_ATOMIC_lane0;
  wire                execute_ctrl3_down_AguPlugin_LOAD_lane0;
  wire                execute_ctrl3_down_MulPlugin_HIGH_lane0;
  wire       [1:0]    execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl3_down_COMPLETION_AT_4_lane0;
  wire                execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl3_down_CfuPlugin_logic_CFU_ENABLE_lane0;
  wire                execute_ctrl3_down_early0_MulPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl3_down_integer_RS2_lane0;
  wire       [1:0]    execute_ctrl3_down_AguPlugin_SIZE_lane0;
  reg                 execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0;
  reg                 execute_ctrl4_up_MMU_HAZARD_lane0;
  reg                 execute_ctrl4_up_MMU_REFILL_lane0;
  reg                 execute_ctrl4_up_MMU_ACCESS_FAULT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  reg                 execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  reg        [31:0]   execute_ctrl4_up_MMU_TRANSLATED_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0;
  reg        [3:0]    execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  reg        [19:0]   execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  reg        [19:0]   execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded;
  reg        [19:0]   execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded;
  reg        [19:0]   execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address;
  reg                 execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault;
  reg        [31:0]   execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  reg        [31:0]   execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  reg        [31:0]   execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  reg        [31:0]   execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_2;
  reg        [31:0]   execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_3;
  reg        [3:0]    execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  reg        [4:0]    execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  reg        [62:0]   execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  reg        [0:0]    execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  reg        [1:0]    execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_1;
  reg        [3:0]    execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0;
  reg        [11:0]   execute_ctrl4_up_Decode_STORE_ID_lane0;
  reg                 execute_ctrl4_up_LsuL1_FLUSH_lane0;
  reg                 execute_ctrl4_up_LsuL1_PREFETCH_lane0;
  reg                 execute_ctrl4_up_LsuL1_INVALID_lane0;
  reg                 execute_ctrl4_up_LsuL1_CLEAN_lane0;
  reg                 execute_ctrl4_up_LsuL1_STORE_lane0;
  reg                 execute_ctrl4_up_LsuL1_ATOMIC_lane0;
  reg                 execute_ctrl4_up_LsuL1_LOAD_lane0;
  reg        [1:0]    execute_ctrl4_up_LsuL1_SIZE_lane0;
  reg        [3:0]    execute_ctrl4_up_LsuL1_MASK_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg        [3:0]    execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  reg        [31:0]   execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  reg        [31:0]   execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0;
  reg        [29:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  reg        [46:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  reg        [46:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  reg        [33:0]   execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 execute_ctrl4_up_AguPlugin_FLOAT_lane0;
  reg                 execute_ctrl4_up_AguPlugin_ATOMIC_lane0;
  reg                 execute_ctrl4_up_AguPlugin_STORE_lane0;
  reg                 execute_ctrl4_up_AguPlugin_LOAD_lane0;
  reg                 execute_ctrl4_up_MulPlugin_HIGH_lane0;
  reg        [1:0]    execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl4_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl4_up_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl4_up_AguPlugin_SEL_lane0;
  reg                 execute_ctrl4_up_CfuPlugin_logic_CFU_ENABLE_lane0;
  reg                 execute_ctrl4_up_early0_MulPlugin_SEL_lane0;
  reg        [1:0]    execute_ctrl4_up_AguPlugin_SIZE_lane0;
  reg        [4:0]    execute_ctrl4_up_RD_PHYS_lane0;
  reg        [15:0]   execute_ctrl4_up_Decode_UOP_ID_lane0;
  reg        [31:0]   execute_ctrl4_up_PC_lane0;
  reg        [11:0]   execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [31:0]   execute_ctrl4_up_Decode_UOP_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl2_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl2_down_MulPlugin_HIGH_lane0;
  wire       [1:0]    execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_4_lane0;
  wire                execute_ctrl2_down_COMPLETION_AT_3_lane0;
  wire                execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0;
  wire                execute_ctrl2_down_early0_MulPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_integer_RS2_lane0;
  wire       [11:0]   execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire                execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0;
  reg        [0:0]    execute_ctrl3_up_MMU_L1_HITS_PRE_VALID_lane0;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_valid;
  reg        [4:0]    execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_virtualAddress;
  reg        [9:0]    execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowRead;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowWrite;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowExecute;
  reg                 execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowUser;
  reg        [2:0]    execute_ctrl3_up_MMU_L0_HITS_PRE_VALID_lane0;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_valid;
  reg        [14:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_virtualAddress;
  reg        [19:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowRead;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowWrite;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowExecute;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowUser;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_valid;
  reg        [14:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_virtualAddress;
  reg        [19:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowRead;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowWrite;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowExecute;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowUser;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_valid;
  reg        [14:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_virtualAddress;
  reg        [19:0]   execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowRead;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowWrite;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowExecute;
  reg                 execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowUser;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0;
  reg        [11:0]   execute_ctrl3_up_Decode_STORE_ID_lane0;
  reg                 execute_ctrl3_up_LsuL1_FLUSH_lane0;
  reg                 execute_ctrl3_up_LsuL1_PREFETCH_lane0;
  reg                 execute_ctrl3_up_LsuL1_INVALID_lane0;
  reg                 execute_ctrl3_up_LsuL1_CLEAN_lane0;
  reg                 execute_ctrl3_up_LsuL1_STORE_lane0;
  reg                 execute_ctrl3_up_LsuL1_ATOMIC_lane0;
  reg                 execute_ctrl3_up_LsuL1_LOAD_lane0;
  reg        [1:0]    execute_ctrl3_up_LsuL1_SIZE_lane0;
  reg        [3:0]    execute_ctrl3_up_LsuL1_MASK_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  reg        [3:0]    execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  reg        [31:0]   execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  reg        [0:0]    execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  reg        [1:0]    execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_1;
  reg        [3:0]    execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  reg                 execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  reg        [31:0]   execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  reg                 execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  reg        [3:0]    execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0;
  reg        [31:0]   execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0;
  reg                 execute_ctrl3_up_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  reg                 execute_ctrl3_up_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  reg                 execute_ctrl3_up_early0_BranchPlugin_logic_alu_EQ_lane0;
  reg        [31:0]   execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  reg        [31:0]   execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  reg        [31:0]   execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  reg        [31:0]   execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0;
  reg        [29:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  reg        [46:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  reg        [46:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  reg        [33:0]   execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  reg                 execute_ctrl3_up_early0_SrcPlugin_LESS_lane0;
  reg        [31:0]   execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 execute_ctrl3_up_AguPlugin_FLOAT_lane0;
  reg                 execute_ctrl3_up_AguPlugin_ATOMIC_lane0;
  reg                 execute_ctrl3_up_AguPlugin_STORE_lane0;
  reg                 execute_ctrl3_up_AguPlugin_LOAD_lane0;
  reg                 execute_ctrl3_up_MulPlugin_HIGH_lane0;
  reg        [1:0]    execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0;
  reg        [1:0]    execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl3_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl3_up_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl3_up_AguPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_CsrAccessPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_CfuPlugin_logic_CFU_ENABLE_lane0;
  reg                 execute_ctrl3_up_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_early0_MulPlugin_SEL_lane0;
  reg                 execute_ctrl3_up_early0_BranchPlugin_SEL_lane0;
  reg        [31:0]   execute_ctrl3_up_integer_RS2_lane0;
  reg        [1:0]    execute_ctrl3_up_AguPlugin_SIZE_lane0;
  reg        [4:0]    execute_ctrl3_up_RD_PHYS_lane0;
  reg        [15:0]   execute_ctrl3_up_Decode_UOP_ID_lane0;
  reg        [31:0]   execute_ctrl3_up_PC_lane0;
  reg        [11:0]   execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg                 execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   execute_ctrl3_up_Decode_UOP_lane0;
  wire       [1:0]    execute_ctrl1_down_AguPlugin_SIZE_lane0;
  wire                execute_ctrl1_down_COMPLETED_lane0;
  wire       [4:0]    execute_ctrl1_down_RD_PHYS_lane0;
  wire       [15:0]   execute_ctrl1_down_Decode_UOP_ID_lane0;
  wire       [11:0]   execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [31:0]   execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0;
  wire                execute_ctrl1_down_isReady;
  reg        [2:0]    execute_ctrl2_up_early0_EnvPlugin_OP_lane0;
  reg                 execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  reg                 execute_ctrl2_up_AguPlugin_FLOAT_lane0;
  reg                 execute_ctrl2_up_AguPlugin_ATOMIC_lane0;
  reg                 execute_ctrl2_up_AguPlugin_STORE_lane0;
  reg                 execute_ctrl2_up_AguPlugin_LOAD_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0;
  reg                 execute_ctrl2_up_DivPlugin_REM_lane0;
  reg                 execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0;
  reg                 execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0;
  reg                 execute_ctrl2_up_MulPlugin_HIGH_lane0;
  reg        [0:0]    execute_ctrl2_up_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0;
  reg        [0:0]    execute_ctrl2_up_CfuPlugin_logic_CFU_ENCODING_lane0;
  reg        [1:0]    execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0;
  reg                 execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0;
  reg                 execute_ctrl2_up_SrcStageables_UNSIGNED_lane0;
  reg                 execute_ctrl2_up_BYPASSED_AT_3_lane0;
  reg        [1:0]    execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  reg                 execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl2_up_SrcStageables_ZERO_lane0;
  reg                 execute_ctrl2_up_SrcStageables_REVERT_lane0;
  reg        [1:0]    execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  reg                 execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0;
  reg                 execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl2_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl2_up_COMPLETION_AT_2_lane0;
  reg                 execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl2_up_AguPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_CsrAccessPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_CfuPlugin_logic_CFU_ENABLE_lane0;
  reg                 execute_ctrl2_up_early0_EnvPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_MulPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0;
  reg                 execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0;
  reg        [31:0]   execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0;
  reg        [1:0]    execute_ctrl2_up_AguPlugin_SIZE_lane0;
  reg        [15:0]   execute_ctrl2_up_Decode_UOP_ID_lane0;
  reg        [31:0]   execute_ctrl2_up_PC_lane0;
  reg        [11:0]   execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [31:0]   execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   execute_ctrl2_up_Decode_UOP_lane0;
  wire                execute_ctrl0_down_COMPLETED_lane0;
  wire       [4:0]    execute_ctrl0_down_RD_PHYS_lane0;
  wire                execute_ctrl0_down_TRAP_lane0;
  wire       [31:0]   execute_ctrl0_down_PC_lane0;
  wire       [11:0]   execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [31:0]   execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0;
  reg        [1:0]    execute_ctrl1_up_AguPlugin_SIZE_lane0;
  reg                 execute_ctrl1_up_COMPLETED_lane0;
  reg        [4:0]    execute_ctrl1_up_RS2_PHYS_lane0;
  reg        [4:0]    execute_ctrl1_up_RS1_PHYS_lane0;
  reg        [15:0]   execute_ctrl1_up_Decode_UOP_ID_lane0;
  reg                 execute_ctrl1_up_TRAP_lane0;
  reg        [31:0]   execute_ctrl1_up_PC_lane0;
  reg        [11:0]   execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0;
  reg        [1:0]    execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  reg        [31:0]   execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  reg                 execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0;
  reg        [31:0]   execute_ctrl1_up_Decode_UOP_lane0;
  wire                decode_ctrls_1_down_isReady;
  wire                decode_ctrls_0_down_Prediction_ALIGN_REDO_0;
  wire       [0:0]    decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [0:0]    decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [31:0]   decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0;
  wire                decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0;
  wire       [11:0]   decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [31:0]   decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0;
  wire                decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0;
  wire       [31:0]   decode_ctrls_0_down_Decode_INSTRUCTION_0;
  wire                decode_ctrls_0_down_isValid;
  wire                decode_ctrls_0_down_isReady;
  reg                 decode_ctrls_1_up_Prediction_ALIGN_REDO_0;
  reg        [0:0]    decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  reg        [0:0]    decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  reg        [31:0]   decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0;
  reg                 decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0;
  reg        [11:0]   decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0;
  reg        [1:0]    decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0;
  reg        [9:0]    decode_ctrls_1_up_Decode_DOP_ID_0;
  reg        [31:0]   decode_ctrls_1_up_PC_0;
  reg        [31:0]   decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0;
  reg                 decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0;
  reg        [31:0]   decode_ctrls_1_up_Decode_INSTRUCTION_0;
  wire       [9:0]    fetch_logic_ctrls_1_down_Fetch_ID;
  wire                fetch_logic_ctrls_1_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_1_down_isValid;
  wire                fetch_logic_ctrls_1_down_isReady;
  reg                 fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT;
  reg                 fetch_logic_ctrls_2_up_MMU_PAGE_FAULT;
  reg                 fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE;
  reg        [31:0]   fetch_logic_ctrls_2_up_MMU_TRANSLATED;
  reg                 fetch_logic_ctrls_2_up_MMU_REFILL;
  reg                 fetch_logic_ctrls_2_up_MMU_HAZARD;
  reg        [0:0]    fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_TAKEN;
  reg        [0:0]    fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_BRANCH;
  reg        [31:0]   fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_PC;
  reg                 fetch_logic_ctrls_2_up_Prediction_WORD_JUMPED;
  reg        [1:0]    fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT;
  reg                 fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_2;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_3;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD;
  reg        [31:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0;
  reg        [31:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1;
  reg        [31:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_2;
  reg        [31:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_3;
  reg        [0:0]    fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  reg        [1:0]    fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_1;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_2_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_2_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_2_address;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_3_loaded;
  reg                 fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_3_error;
  reg        [19:0]   fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_3_address;
  reg        [11:0]   fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY;
  reg        [9:0]    fetch_logic_ctrls_2_up_Fetch_ID;
  reg                 fetch_logic_ctrls_2_up_Fetch_PC_FAULT;
  reg        [31:0]   fetch_logic_ctrls_2_up_Fetch_WORD_PC;
  wire                fetch_logic_ctrls_0_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_0_down_isValid;
  reg        [0:0]    fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS;
  reg                 fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid;
  reg        [13:0]   fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address;
  reg        [1:0]    fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0;
  reg        [11:0]   fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY;
  reg        [13:0]   fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH;
  reg        [5:0]    fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  reg        [0:0]    fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  reg        [1:0]    fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_1;
  reg                 fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg                 _zz_1;
  reg        [9:0]    fetch_logic_ctrls_1_up_Fetch_ID;
  reg                 fetch_logic_ctrls_1_up_Fetch_PC_FAULT;
  reg        [31:0]   fetch_logic_ctrls_1_up_Fetch_WORD_PC;
  reg                 fetch_logic_ctrls_2_up_valid;
  wire                decode_ctrls_1_down_valid;
  reg                 fetch_logic_ctrls_1_down_valid;
  wire                decode_ctrls_0_down_valid;
  reg                 fetch_logic_ctrls_0_down_valid;
  wire                execute_ctrl0_up_ready;
  wire                execute_ctrl0_down_ready;
  wire                execute_ctrl1_up_ready;
  wire                execute_ctrl1_down_ready;
  wire                execute_ctrl2_up_ready;
  wire                execute_ctrl2_down_ready;
  wire                execute_ctrl3_up_ready;
  wire                execute_ctrl3_down_ready;
  wire                fetch_logic_ctrls_0_down_ready;
  wire                execute_ctrl4_up_ready;
  wire                decode_ctrls_0_up_ready;
  wire                fetch_logic_ctrls_1_up_cancel;
  wire                execute_ctrl4_down_ready;
  reg                 decode_ctrls_0_down_ready;
  wire                fetch_logic_ctrls_1_down_ready;
  wire                execute_ctrl5_up_ready;
  wire                fetch_logic_ctrls_2_up_ready;
  wire                fetch_logic_ctrls_2_up_cancel;
  wire                execute_ctrl5_down_ready;
  wire                execute_ctrl4_down_AguPlugin_ATOMIC_lane0;
  wire       [11:0]   execute_ctrl4_down_Decode_STORE_ID_lane0;
  wire       [31:0]   execute_ctrl4_down_MMU_TRANSLATED_lane0;
  wire       [1:0]    execute_ctrl4_down_AguPlugin_SIZE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl4_down_AguPlugin_LOAD_lane0;
  wire                execute_ctrl4_down_RD_ENABLE_lane0;
  reg                 execute_ctrl4_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl4_LANE_SEL_lane0_bypass;
  wire                execute_ctrl3_down_RD_ENABLE_lane0;
  reg                 execute_ctrl3_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl3_LANE_SEL_lane0_bypass;
  wire                execute_ctrl2_down_RD_ENABLE_lane0;
  reg                 execute_ctrl2_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl2_LANE_SEL_lane0_bypass;
  wire                execute_ctrl1_down_RD_ENABLE_lane0;
  reg                 execute_ctrl1_RD_ENABLE_lane0_bypass;
  wire                execute_ctrl1_down_LANE_SEL_lane0;
  reg                 execute_ctrl1_LANE_SEL_lane0_bypass;
  wire                execute_ctrl0_down_RD_ENABLE_lane0;
  reg                 execute_ctrl0_RD_ENABLE_lane0_bypass;
  reg                 execute_ctrl0_LANE_SEL_lane0_bypass;
  wire                execute_ctrl1_down_TRAP_lane0;
  wire       [2:0]    execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
  wire                execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
  wire                execute_ctrl1_down_AguPlugin_INVALIDATE_lane0;
  wire                execute_ctrl1_down_AguPlugin_CLEAN_lane0;
  wire                execute_ctrl1_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
  wire                execute_ctrl1_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl1_down_AguPlugin_LOAD_lane0;
  wire                execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire                execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire                execute_ctrl1_down_DivPlugin_REM_lane0;
  wire                execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire                execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire                execute_ctrl1_down_MulPlugin_HIGH_lane0;
  wire       [0:0]    execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0;
  wire       [0:0]    execute_ctrl1_down_CfuPlugin_logic_CFU_ENCODING_lane0;
  wire       [1:0]    execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
  wire                execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_3_lane0;
  wire       [1:0]    execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  wire                execute_ctrl1_down_SrcStageables_ZERO_lane0;
  wire                execute_ctrl1_down_SrcStageables_REVERT_lane0;
  wire       [1:0]    execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  reg                 execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl1_down_COMPLETION_AT_2_lane0;
  reg                 execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
  reg                 execute_ctrl1_down_AguPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0;
  reg                 execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
  reg                 execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
  wire                execute_ctrl4_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                execute_ctrl3_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                execute_ctrl2_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  wire       [4:0]    execute_ctrl1_down_RS2_PHYS_lane0;
  wire       [4:0]    execute_ctrl0_down_RS2_PHYS_lane0;
  wire       [31:0]   execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [4:0]    execute_ctrl5_down_RD_PHYS_lane0;
  reg                 execute_ctrl5_up_RD_ENABLE_lane0;
  reg                 execute_ctrl5_up_LANE_SEL_lane0;
  wire       [4:0]    execute_ctrl3_down_RD_PHYS_lane0;
  wire       [4:0]    execute_ctrl1_down_RS1_PHYS_lane0;
  wire       [4:0]    execute_ctrl0_down_RS1_PHYS_lane0;
  reg                 _zz_2;
  wire                execute_ctrl3_down_CsrAccessPlugin_SEL_lane0;
  wire       [4:0]    execute_ctrl2_down_RD_PHYS_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0;
  wire                execute_ctrl2_down_CsrAccessPlugin_SEL_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT;
  reg                 fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT;
  reg                 fetch_logic_ctrls_1_down_MMU_PAGE_FAULT;
  reg                 fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE;
  reg                 fetch_logic_ctrls_1_down_MMU_ALLOW_READ;
  reg                 fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE;
  reg        [31:0]   fetch_logic_ctrls_1_down_MMU_TRANSLATED;
  reg                 fetch_logic_ctrls_1_down_MMU_REFILL;
  reg                 fetch_logic_ctrls_1_down_MMU_HAZARD;
  wire       [0:0]    fetch_logic_ctrls_1_down_MMU_L1_HITS;
  wire       [0:0]    fetch_logic_ctrls_1_down_MMU_L1_HITS_PRE_VALID;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid;
  wire       [4:0]    fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_virtualAddress;
  wire       [9:0]    fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowRead;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowWrite;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowExecute;
  wire                fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowUser;
  reg        [1:0]    fetch_logic_ctrls_1_down_MMU_L0_HITS;
  reg        [1:0]    fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid;
  wire       [14:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_virtualAddress;
  wire       [19:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowRead;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowWrite;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowExecute;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowUser;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid;
  wire       [14:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_virtualAddress;
  wire       [19:0]   fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowRead;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowWrite;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowExecute;
  wire                fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowUser;
  wire       [31:0]   execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_0;
  wire       [31:0]   execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_1;
  wire       [31:0]   execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_2;
  wire       [31:0]   execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_3;
  wire       [3:0]    execute_ctrl3_down_MMU_WAYS_OH_lane0;
  wire                execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0;
  reg                 execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid;
  wire       [4:0]    execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_virtualAddress;
  wire       [9:0]    execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowRead;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowWrite;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowExecute;
  wire                execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowUser;
  wire       [0:0]    execute_ctrl3_down_MMU_L1_HITS_PRE_VALID_lane0;
  wire       [0:0]    execute_ctrl3_down_MMU_L1_HITS_lane0;
  wire       [0:0]    execute_ctrl2_down_MMU_L1_HITS_PRE_VALID_lane0;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid;
  wire       [4:0]    execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_virtualAddress;
  wire       [9:0]    execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowRead;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowWrite;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowExecute;
  wire                execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowUser;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid;
  wire       [14:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_virtualAddress;
  wire       [19:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowRead;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowWrite;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowExecute;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowUser;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid;
  wire       [14:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_virtualAddress;
  wire       [19:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowRead;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowWrite;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowExecute;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowUser;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_valid;
  wire       [14:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_virtualAddress;
  wire       [19:0]   execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowRead;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowWrite;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowExecute;
  wire                execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowUser;
  wire       [2:0]    execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0;
  reg        [2:0]    execute_ctrl3_down_MMU_L0_HITS_lane0;
  reg        [2:0]    execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid;
  wire       [14:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_virtualAddress;
  wire       [19:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowRead;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowWrite;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowExecute;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowUser;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid;
  wire       [14:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_virtualAddress;
  wire       [19:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowRead;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowWrite;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowExecute;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowUser;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid;
  wire       [14:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_virtualAddress;
  wire       [19:0]   execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowRead;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowWrite;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowExecute;
  wire                execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowUser;
  wire                fetch_logic_ctrls_0_up_isFiring;
  reg        [9:0]    fetch_logic_ctrls_0_up_Fetch_ID;
  wire                fetch_logic_ctrls_0_up_Fetch_PC_FAULT;
  wire       [31:0]   fetch_logic_ctrls_0_up_Fetch_WORD_PC;
  reg                 fetch_logic_ctrls_0_up_ready;
  wire                fetch_logic_ctrls_0_up_valid;
  reg                 PcPlugin_logic_harts_0_aggregator_fault_1;
  reg        [31:0]   PcPlugin_logic_harts_0_aggregator_target_1;
  wire                execute_ctrl4_down_AguPlugin_FLOAT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 execute_ctrl4_up_COMMIT_lane0;
  reg                 execute_ctrl4_COMMIT_lane0_bypass;
  reg                 execute_ctrl4_up_TRAP_lane0;
  reg                 execute_ctrl4_TRAP_lane0_bypass;
  wire                execute_ctrl4_down_AguPlugin_SEL_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  wire                execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0;
  wire                execute_ctrl4_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  wire                execute_ctrl4_down_MMU_HAZARD_lane0;
  wire                execute_ctrl4_down_MMU_REFILL_lane0;
  wire                execute_ctrl4_down_MMU_ACCESS_FAULT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  wire                execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  wire                execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  wire       [31:0]   execute_ctrl4_down_integer_RS2_lane0;
  wire       [31:0]   execute_ctrl4_down_Decode_UOP_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1_SIZE_lane0;
  wire                execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0;
  reg        [31:0]   execute_ctrl4_up_integer_RS2_lane0;
  reg                 execute_ctrl3_down_MMU_HAZARD_lane0;
  reg                 execute_ctrl3_down_MMU_REFILL_lane0;
  reg                 execute_ctrl3_down_MMU_ACCESS_FAULT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0;
  reg                 execute_ctrl3_down_MMU_ALLOW_READ_lane0;
  reg                 execute_ctrl3_down_MMU_ALLOW_WRITE_lane0;
  wire                execute_ctrl3_down_AguPlugin_STORE_lane0;
  reg                 execute_ctrl3_down_MMU_PAGE_FAULT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  wire       [31:0]   execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  reg                 execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  wire                execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  wire                execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  wire                execute_ctrl3_down_LsuL1_ATOMIC_lane0;
  wire                execute_ctrl3_down_AguPlugin_SEL_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  reg                 execute_ctrl4_LsuL1_SEL_lane0_bypass;
  wire                execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0;
  reg                 execute_ctrl4_up_LsuL1_SEL_lane0;
  reg                 execute_ctrl3_LsuL1_SEL_lane0_bypass;
  wire                execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0;
  reg                 execute_ctrl3_up_LsuL1_SEL_lane0;
  reg        [31:0]   execute_ctrl3_down_MMU_TRANSLATED_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0;
  wire       [11:0]   execute_ctrl2_down_Decode_STORE_ID_lane0;
  wire                execute_ctrl2_down_LsuL1_FLUSH_lane0;
  wire                execute_ctrl2_down_LsuL1_PREFETCH_lane0;
  wire                execute_ctrl2_down_LsuL1_INVALID_lane0;
  wire                execute_ctrl2_down_LsuL1_CLEAN_lane0;
  wire                execute_ctrl2_down_LsuL1_STORE_lane0;
  wire                execute_ctrl2_down_LsuL1_ATOMIC_lane0;
  wire                execute_ctrl2_down_LsuL1_LOAD_lane0;
  wire       [1:0]    execute_ctrl2_down_LsuL1_SIZE_lane0;
  wire       [3:0]    execute_ctrl2_down_LsuL1_MASK_lane0;
  wire                execute_ctrl2_down_LsuL1_SEL_lane0;
  wire                execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
  wire                execute_ctrl2_down_AguPlugin_STORE_lane0;
  wire                execute_ctrl2_down_AguPlugin_LOAD_lane0;
  wire       [1:0]    execute_ctrl2_down_AguPlugin_SIZE_lane0;
  wire                execute_ctrl2_down_AguPlugin_SEL_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0;
  wire                execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  wire                execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0;
  wire       [1:0]    execute_ctrl3_down_LsuL1_SIZE_lane0;
  wire                execute_ctrl3_down_LsuL1_STORE_lane0;
  wire                execute_ctrl3_down_LsuL1_LOAD_lane0;
  wire       [11:0]   execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [31:0]   execute_ctrl4_down_PC_lane0;
  wire                execute_ctrl4_down_TRAP_lane0;
  wire                execute_ctrl5_down_COMMIT_lane0;
  wire                execute_ctrl5_down_isReady;
  wire                execute_ctrl5_down_LANE_SEL_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1_READ_DATA_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire       [3:0]    execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire       [3:0]    execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  reg        [31:0]   execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0;
  wire       [3:0]    execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  wire       [31:0]   execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  wire                execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0;
  wire       [3:0]    execute_ctrl4_down_LsuL1_MASK_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  wire       [0:0]    execute_ctrl4_down_LsuL1_WAIT_WRITEBACK_lane0;
  wire       [0:0]    execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
  wire                execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0;
  wire                execute_ctrl4_down_LsuL1_INVALID_lane0;
  wire                execute_ctrl4_down_LsuL1_CLEAN_lane0;
  wire                execute_ctrl4_up_isReady;
  wire                execute_ctrl4_down_LsuL1_REFILL_HIT_lane0;
  wire                execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0;
  wire                execute_ctrl4_down_LsuL1_FAULT_lane0;
  wire                execute_ctrl4_down_LsuL1_MISS_lane0;
  wire                execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0;
  wire                execute_ctrl4_down_LsuL1_HAZARD_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0;
  wire                execute_ctrl4_down_LsuL1_ABORD_lane0;
  wire                execute_ctrl4_down_LsuL1_PREFETCH_lane0;
  wire                execute_ctrl4_down_LsuL1_LOAD_lane0;
  wire       [3:0]    execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  wire       [19:0]   execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  wire       [19:0]   execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded;
  wire       [19:0]   execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded;
  wire       [19:0]   execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault;
  wire       [0:0]    execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  wire       [1:0]    execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_1;
  wire       [3:0]    execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire                execute_ctrl4_down_LsuL1_ATOMIC_lane0;
  wire                execute_ctrl4_down_LsuL1_STORE_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0;
  wire                execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0;
  reg        [3:0]    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
  wire       [0:0]    execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  wire       [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_1;
  wire       [3:0]    execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire       [0:0]    execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0;
  wire       [1:0]    execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_1;
  wire       [3:0]    execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty;
  wire       [0:0]    execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  wire       [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_1;
  wire       [3:0]    execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  wire       [19:0]   execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  wire       [19:0]   execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded;
  wire       [19:0]   execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded;
  wire       [19:0]   execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault;
  reg        [0:0]    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  reg        [1:0]    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_1;
  reg        [3:0]    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  wire       [0:0]    execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  wire       [1:0]    execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_1;
  wire       [3:0]    execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  wire                execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  wire                execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  wire       [31:0]   execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  wire                execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  reg        [1:0]    execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [31:0]   execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [31:0]   execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2;
  wire       [31:0]   execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3;
  wire       [3:0]    execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
  wire       [31:0]   execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
  wire       [31:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  wire       [31:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  wire       [31:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2;
  wire       [31:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3;
  wire       [3:0]    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
  reg        [3:0]    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_2;
  wire       [63:0]   execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_3;
  reg        [3:0]    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
  wire       [31:0]   execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0;
  reg                 _zz_3;
  reg                 _zz_4;
  wire                decode_ctrls_0_down_TRAP_0;
  wire                decode_ctrls_1_down_LANE_SEL_0;
  reg                 decode_ctrls_1_LANE_SEL_0_bypass;
  wire                decode_ctrls_0_down_LANE_SEL_0;
  reg                 decode_ctrls_0_LANE_SEL_0_bypass;
  wire                decode_ctrls_0_up_isMoving;
  wire       [31:0]   fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC;
  wire       [0:0]    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN;
  wire       [0:0]    fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH;
  wire       [11:0]   fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY;
  wire       [1:0]    fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0;
  wire       [9:0]    fetch_logic_ctrls_2_down_Fetch_ID;
  wire                fetch_logic_ctrls_2_down_ready;
  wire                fetch_logic_ctrls_2_down_valid;
  wire                fetch_logic_ctrls_2_down_isValid;
  wire       [0:0]    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN;
  wire       [0:0]    fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH;
  wire       [11:0]   fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
  wire       [31:0]   fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_PC;
  wire                fetch_logic_ctrls_1_down_Prediction_WORD_JUMPED;
  wire                fetch_logic_ctrls_1_up_isCancel;
  wire                fetch_logic_ctrls_1_up_isReady;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
  wire       [0:0]    fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS;
  wire                fetch_logic_ctrls_1_up_isValid;
  wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT;
  (* keep , syn_keep *) wire       [15:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [29:0]   fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop /* synthesis syn_keep = 1 */ ;
  wire       [0:0]    fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS;
  wire       [15:0]   execute_ctrl0_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl0_down_isReady;
  wire                execute_ctrl0_down_LANE_SEL_lane0;
  wire       [9:0]    decode_ctrls_1_down_Decode_DOP_ID_0;
  wire                decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0;
  wire                decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0;
  wire       [4:0]    execute_ctrl4_down_RD_PHYS_lane0;
  wire                execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire       [15:0]   execute_ctrl4_down_Decode_UOP_ID_lane0;
  wire                execute_ctrl4_down_COMMIT_lane0;
  reg                 execute_ctrl4_up_RD_ENABLE_lane0;
  wire                execute_ctrl4_down_LANE_SEL_lane0;
  wire       [31:0]   execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [31:0]   execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  reg                 execute_ctrl3_up_RD_ENABLE_lane0;
  wire                execute_ctrl3_down_LANE_SEL_lane0;
  wire       [31:0]   execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  reg        [31:0]   execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire                execute_ctrl2_down_LANE_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  wire       [31:0]   execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  wire                execute_ctrl0_up_COMPLETED_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0;
  wire       [4:0]    execute_ctrl0_up_RD_PHYS_lane0;
  reg                 execute_ctrl0_up_RD_ENABLE_lane0;
  wire       [4:0]    execute_ctrl0_up_RS2_PHYS_lane0;
  wire                execute_ctrl0_up_RS2_ENABLE_lane0;
  wire       [4:0]    execute_ctrl0_up_RS1_PHYS_lane0;
  wire                execute_ctrl0_up_RS1_ENABLE_lane0;
  wire       [15:0]   execute_ctrl0_up_Decode_UOP_ID_lane0;
  wire                execute_ctrl0_up_TRAP_lane0;
  wire       [31:0]   execute_ctrl0_up_PC_lane0;
  wire                execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0;
  wire                execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0;
  reg                 execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0;
  wire                execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0;
  wire       [11:0]   execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0;
  wire       [1:0]    execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [0:0]    execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0;
  wire       [0:0]    execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0;
  wire       [31:0]   execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  wire       [31:0]   execute_ctrl0_up_Decode_UOP_lane0;
  wire                execute_ctrl0_up_LANE_SEL_lane0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  wire                decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  wire                decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  wire                decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  wire                decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  wire                decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  wire                decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  wire       [11:0]   decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [0:0]    decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [0:0]    decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [31:0]   decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0;
  wire                decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
  wire                decode_ctrls_1_up_isValid;
  reg                 decode_ctrls_1_down_ready;
  wire                execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0;
  wire                execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0;
  wire                execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
  wire                execute_ctrl2_down_BYPASSED_AT_3_lane0;
  reg        [4:0]    execute_ctrl2_up_RD_PHYS_lane0;
  reg                 execute_ctrl2_up_RD_ENABLE_lane0;
  wire                execute_ctrl1_down_BYPASSED_AT_2_lane0;
  reg        [4:0]    execute_ctrl1_up_RD_PHYS_lane0;
  reg                 execute_ctrl1_up_RD_ENABLE_lane0;
  wire       [31:0]   decode_ctrls_1_down_Decode_UOP_0;
  reg                 decode_ctrls_1_up_TRAP_0;
  reg                 decode_ctrls_1_TRAP_0_bypass;
  wire       [15:0]   decode_ctrls_1_down_Decode_UOP_ID_0;
  wire                decode_ctrls_1_up_isReady;
  wire                decode_ctrls_1_down_TRAP_0;
  wire       [31:0]   decode_ctrls_1_down_PC_0;
  wire                decode_ctrls_1_down_Prediction_ALIGN_REDO_0;
  wire                decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0;
  reg                 decode_ctrls_1_up_LANE_SEL_0;
  wire       [31:0]   decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0;
  wire                decode_ctrls_1_down_CfuPlugin_logic_CFU_ENABLE_0;
  wire                decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0;
  reg                 decode_ctrls_1_down_Decode_LEGAL_0;
  wire       [4:0]    decode_ctrls_1_down_RD_PHYS_0;
  reg                 decode_ctrls_1_down_RD_ENABLE_0;
  wire       [4:0]    decode_ctrls_1_down_RS2_PHYS_0;
  wire                decode_ctrls_1_down_RS2_ENABLE_0;
  wire       [4:0]    decode_ctrls_1_down_RS1_PHYS_0;
  wire       [31:0]   decode_ctrls_1_down_Decode_INSTRUCTION_0;
  wire                decode_ctrls_1_down_RS1_ENABLE_0;
  wire                decode_ctrls_1_up_isCanceling;
  wire                decode_ctrls_1_up_ready;
  reg                 decode_ctrls_1_up_valid;
  wire                decode_ctrls_1_up_isMoving;
  wire                execute_ctrl4_down_COMPLETION_AT_4_lane0;
  reg                 execute_ctrl4_up_COMPLETED_lane0;
  wire                execute_ctrl4_down_COMPLETED_lane0;
  wire                execute_ctrl4_COMPLETED_lane0_bypass;
  wire                execute_ctrl3_down_COMPLETION_AT_3_lane0;
  reg                 execute_ctrl3_up_COMPLETED_lane0;
  wire                execute_ctrl3_down_COMPLETED_lane0;
  wire                execute_ctrl3_COMPLETED_lane0_bypass;
  wire                execute_ctrl2_down_COMPLETION_AT_2_lane0;
  reg                 execute_ctrl2_up_COMPLETED_lane0;
  wire                execute_ctrl2_down_COMPLETED_lane0;
  wire                execute_ctrl2_COMPLETED_lane0_bypass;
  reg                 execute_ctrl1_up_LANE_SEL_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
  wire       [1:0]    execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  wire       [31:0]   execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  wire                execute_ctrl3_down_isReady;
  wire                execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0;
  wire                execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0;
  reg                 execute_ctrl3_up_COMMIT_lane0;
  wire                execute_ctrl3_down_COMMIT_lane0;
  reg                 execute_ctrl3_COMMIT_lane0_bypass;
  reg                 execute_ctrl3_up_TRAP_lane0;
  wire                execute_ctrl3_down_TRAP_lane0;
  reg                 execute_ctrl3_TRAP_lane0_bypass;
  wire                execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0;
  wire       [15:0]   execute_ctrl3_down_Decode_UOP_ID_lane0;
  reg        [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter_1;
  wire       [11:0]   execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
  wire       [31:0]   execute_ctrl3_down_PC_lane0;
  wire                execute_ctrl3_down_early0_BranchPlugin_SEL_lane0;
  wire                execute_ctrl3_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire                execute_ctrl3_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  wire                execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0;
  wire       [31:0]   execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  wire       [31:0]   execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  wire       [31:0]   execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  wire                execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  wire                execute_ctrl3_down_early0_SrcPlugin_LESS_lane0;
  wire                execute_ctrl3_down_early0_BranchPlugin_logic_alu_EQ_lane0;
  wire       [31:0]   execute_ctrl3_down_Decode_UOP_lane0;
  wire       [1:0]    execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  wire       [31:0]   execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0;
  wire                execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0;
  wire                execute_ctrl2_up_COMMIT_lane0;
  wire                execute_ctrl2_down_COMMIT_lane0;
  reg                 execute_ctrl2_COMMIT_lane0_bypass;
  reg                 execute_ctrl2_up_TRAP_lane0;
  wire                execute_ctrl2_down_TRAP_lane0;
  reg                 execute_ctrl2_TRAP_lane0_bypass;
  wire                execute_ctrl2_down_early0_EnvPlugin_SEL_lane0;
  wire                execute_ctrl4_down_LsuL1_FLUSH_lane0;
  wire                execute_ctrl4_down_LsuL1_SEL_lane0;
  wire                execute_ctrl3_down_LsuL1_FLUSH_lane0;
  wire                execute_ctrl3_down_LsuL1_SEL_lane0;
  wire       [31:0]   execute_ctrl0_down_Decode_UOP_lane0;
  reg                 execute_ctrl4_up_CfuPlugin_logic_CFU_IN_FLIGHT_lane0;
  reg                 execute_ctrl3_up_CfuPlugin_logic_CFU_IN_FLIGHT_lane0;
  wire                execute_ctrl4_down_isReady;
  wire                execute_ctrl4_down_CfuPlugin_logic_CFU_ENABLE_lane0;
  wire                execute_ctrl4_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0;
  wire       [0:0]    execute_ctrl2_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0;
  wire       [0:0]    execute_ctrl2_down_CfuPlugin_logic_CFU_ENCODING_lane0;
  wire                decode_ctrls_0_up_isValid;
  wire                decode_ctrls_0_up_valid;
  wire                decode_ctrls_0_up_Prediction_ALIGN_REDO_0;
  wire       [0:0]    decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  wire       [0:0]    decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  wire       [31:0]   decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0;
  wire                decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0;
  wire                decode_ctrls_0_up_TRAP_0;
  wire                decode_ctrls_0_up_Prediction_WORD_JUMPED_0;
  wire       [31:0]   decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0;
  wire       [0:0]    decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0;
  wire       [0:0]    decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0;
  wire       [11:0]   decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0;
  wire       [1:0]    decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0;
  wire       [9:0]    decode_ctrls_0_up_Fetch_ID_0;
  wire       [9:0]    decode_ctrls_0_up_Decode_DOP_ID_0;
  wire       [31:0]   decode_ctrls_0_up_PC_0;
  reg        [31:0]   decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0;
  wire                decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0;
  wire       [31:0]   decode_ctrls_0_up_Decode_INSTRUCTION_0;
  wire                decode_ctrls_0_up_isFiring;
  wire       [0:0]    fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST;
  wire                fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED;
  wire       [0:0]    fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK;
  (* keep , syn_keep *) wire       [31:0]   execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [31:0]   execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) reg        [31:0]   execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 /* synthesis syn_keep = 1 */ ;
  wire       [1:0]    execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire       [31:0]   execute_ctrl2_down_Decode_UOP_lane0;
  reg                 execute_ctrl3_up_LANE_SEL_lane0;
  wire       [1:0]    execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  wire                execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  reg                 execute_ctrl4_up_LANE_SEL_lane0;
  wire                execute_ctrl2_down_SrcStageables_UNSIGNED_lane0;
  wire                execute_ctrl2_down_SrcStageables_ZERO_lane0;
  wire                execute_ctrl2_down_SrcStageables_REVERT_lane0;
  wire       [31:0]   execute_ctrl1_down_PC_lane0;
  wire       [31:0]   execute_ctrl1_down_integer_RS2_lane0;
  wire       [1:0]    execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0;
  wire       [31:0]   execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   execute_ctrl1_down_integer_RS1_lane0;
  wire       [0:0]    execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0;
  wire       [31:0]   execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  wire       [31:0]   execute_ctrl1_down_Decode_UOP_lane0;
  wire       [2:0]    execute_ctrl2_down_early0_EnvPlugin_OP_lane0;
  wire       [31:0]   execute_ctrl2_down_PC_lane0;
  wire       [15:0]   execute_ctrl2_down_Decode_UOP_ID_lane0;
  wire                decode_ctrls_1_lane0_upIsCancel;
  wire                decode_ctrls_1_lane0_downIsCancel;
  wire       [9:0]    decode_ctrls_0_down_Decode_DOP_ID_0;
  wire       [9:0]    decode_ctrls_0_down_Fetch_ID_0;
  wire       [31:0]   decode_ctrls_0_down_PC_0;
  wire                decode_ctrls_0_up_isReady;
  wire                decode_ctrls_0_up_LANE_SEL_0;
  wire                decode_ctrls_0_lane0_upIsCancel;
  wire                decode_ctrls_0_lane0_downIsCancel;
  wire       [9:0]    fetch_logic_ctrls_0_down_Fetch_ID;
  reg                 _zz_wr_en;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_pop_aheadValue;
  wire       [13:0]   fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH;
  wire                fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid;
  wire       [13:0]   fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0;
  wire                fetch_logic_ctrls_0_down_isReady;
  (* keep , syn_keep *) reg        [1:0]    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 /* synthesis syn_keep = 1 */ ;
  wire                fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid;
  wire       [13:0]   fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address;
  wire       [1:0]    fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0;
  wire       [11:0]   fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
  wire       [13:0]   fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  reg                 _zz_5;
  wire       [1:0]    execute_ctrl0_down_AguPlugin_SIZE_lane0;
  wire                fetch_logic_ctrls_2_up_isMoving;
  wire                fetch_logic_ctrls_2_up_isCanceling;
  wire                fetch_logic_ctrls_2_down_isReady;
  wire                fetch_logic_ctrls_2_down_TRAP;
  wire                fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION;
  wire                fetch_logic_ctrls_2_down_Fetch_PC_FAULT;
  wire                fetch_logic_ctrls_2_down_MMU_HAZARD;
  wire                fetch_logic_ctrls_2_down_MMU_REFILL;
  wire                fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT;
  wire                fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE;
  wire                fetch_logic_ctrls_2_down_MMU_PAGE_FAULT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT;
  wire                fetch_logic_ctrls_2_up_isCancel;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_2_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_2_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_2_address;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_3_loaded;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_3_error;
  wire       [19:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_3_address;
  wire       [31:0]   fetch_logic_ctrls_2_down_Fetch_WORD_PC;
  wire                fetch_logic_ctrls_2_up_isReady;
  wire                fetch_logic_ctrls_2_up_isValid;
  wire       [0:0]    fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  wire       [1:0]    fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_1;
  wire       [31:0]   fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT;
  wire                fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_2;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_3;
  wire       [2:0]    fetch_logic_ctrls_1_down_MMU_WAYS_OH;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1;
  wire       [31:0]   fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2;
  wire       [5:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD;
  wire       [31:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [31:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire       [31:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_2;
  wire       [31:0]   fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_3;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_2;
  wire                fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_3;
  wire       [31:0]   fetch_logic_ctrls_2_down_Fetch_WORD;
  wire       [31:0]   fetch_logic_ctrls_1_down_Fetch_WORD_PC;
  wire       [31:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  wire       [31:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  wire       [31:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2;
  wire       [31:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3;
  wire       [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  wire       [1:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_1;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg        [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  reg        [1:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_1;
  wire       [5:0]    fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  wire       [0:0]    fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  wire       [1:0]    fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_1;
  wire                fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  reg                 fetch_logic_ctrls_1_up_valid;
  wire                fetch_logic_ctrls_1_up_ready;
  wire       [31:0]   fetch_logic_ctrls_0_down_Fetch_WORD_PC;
  reg                 _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217;
  wire       [0:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0;
  wire       [1:0]    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_1;
  reg                 _zz_6;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_address;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_loaded;
  wire                fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_error;
  wire       [19:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_address;
  reg                 _zz_7;
  reg                 _zz_8;
  reg                 _zz_9;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_2;
  wire       [63:0]   fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_3;
  reg                 _zz_10;
  wire                fetch_logic_ctrls_0_down_isFiring;
  wire       [31:0]   execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0;
  wire                execute_ctrl3_down_early0_DivPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
  wire                execute_ctrl2_down_early0_DivPlugin_SEL_lane0;
  wire                execute_ctrl2_down_isReady;
  wire                execute_ctrl2_down_DivPlugin_REM_lane0;
  wire       [31:0]   execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  wire       [31:0]   execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0;
  wire       [31:0]   execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0;
  wire       [31:0]   execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0;
  wire                execute_ctrl4_down_MulPlugin_HIGH_lane0;
  wire                execute_ctrl4_down_early0_MulPlugin_SEL_lane0;
  wire       [65:0]   execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0;
  wire       [4:0]    execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  wire       [62:0]   execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  wire       [29:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [46:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [46:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  wire       [4:0]    execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  wire       [62:0]   execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  wire       [29:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [46:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [46:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  wire       [29:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  wire       [46:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  wire       [46:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  wire       [33:0]   execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire       [32:0]   execute_ctrl2_down_MUL_SRC2_lane0;
  wire                execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
  wire       [32:0]   execute_ctrl2_down_MUL_SRC1_lane0;
  reg        [31:0]   execute_ctrl2_up_integer_RS2_lane0;
  reg        [31:0]   execute_ctrl2_up_integer_RS1_lane0;
  wire                execute_ctrl2_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0;
  wire                execute_ctrl2_down_CfuPlugin_logic_CFU_ENABLE_lane0;
  reg                 execute_ctrl2_up_LANE_SEL_lane0;
  wire                execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  wire                execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0;
  wire                execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0;
  wire                execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0;
  wire                execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0;
  wire                execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
  wire                execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0;
  wire       [31:0]   execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
  wire       [1:0]    execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire                early0_BranchPlugin_logic_events_branchMiss;
  wire                early0_BranchPlugin_logic_events_branchCount;
  reg                 MmuPlugin_api_fetchTranslationEnable;
  reg                 MmuPlugin_api_lsuTranslationEnable;
  wire                AlignerPlugin_api_singleFetch;
  wire                AlignerPlugin_api_downMoving;
  wire                AlignerPlugin_api_haltIt;
  reg                 DispatchPlugin_api_haltDispatch;
  wire                execute_freeze_valid;
  wire       [0:0]    execute_lane0_api_hartsInflight;
  wire                execute_lane0_ctrls_2_upIsCancel;
  wire                execute_lane0_ctrls_2_downIsCancel;
  reg                 CsrRamPlugin_api_holdRead;
  reg                 CsrRamPlugin_api_holdWrite;
  reg                 CsrAccessPlugin_bus_decode_exception;
  wire                CsrAccessPlugin_bus_decode_read;
  wire                CsrAccessPlugin_bus_decode_write;
  wire       [11:0]   CsrAccessPlugin_bus_decode_address;
  reg                 CsrAccessPlugin_bus_decode_trap;
  wire                PrivilegedPlugin_api_lsuTriggerBus_load;
  wire                PrivilegedPlugin_api_lsuTriggerBus_store;
  reg                 TrapPlugin_api_harts_0_redo;
  reg                 TrapPlugin_api_harts_0_askWake;
  reg                 TrapPlugin_api_harts_0_rvTrap;
  wire                TrapPlugin_api_harts_0_fsmBusy;
  reg                 MmuPlugin_logic_accessBus_cmd_valid;
  wire                MmuPlugin_logic_accessBus_cmd_ready;
  wire       [31:0]   MmuPlugin_logic_accessBus_cmd_payload_address;
  wire       [1:0]    MmuPlugin_logic_accessBus_cmd_payload_size;
  wire                MmuPlugin_logic_accessBus_rsp_valid;
  wire       [31:0]   MmuPlugin_logic_accessBus_rsp_payload_data;
  reg                 MmuPlugin_logic_accessBus_rsp_payload_error;
  reg                 MmuPlugin_logic_accessBus_rsp_payload_redo;
  wire                MmuPlugin_logic_accessBus_rsp_payload_waitAny;
  reg        [0:0]    MmuPlugin_logic_satp_mode;
  reg        [19:0]   MmuPlugin_logic_satp_ppn;
  reg                 MmuPlugin_logic_status_mxr;
  reg                 MmuPlugin_logic_status_sum;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2;
  wire                BtbPlugin_logic_pcPort_valid;
  wire                BtbPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   BtbPlugin_logic_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid;
  wire                BtbPlugin_logic_historyPort_valid;
  wire       [11:0]   BtbPlugin_logic_historyPort_payload_history;
  wire                BtbPlugin_logic_flushPort_valid;
  wire                BtbPlugin_logic_flushPort_payload_self;
  wire                FetchL1Plugin_logic_bus_cmd_valid;
  wire                FetchL1Plugin_logic_bus_cmd_ready;
  wire       [31:0]   FetchL1Plugin_logic_bus_cmd_payload_address;
  wire                FetchL1Plugin_logic_bus_cmd_payload_io;
  wire                FetchL1Plugin_logic_bus_rsp_valid;
  wire                FetchL1Plugin_logic_bus_rsp_ready;
  wire       [63:0]   FetchL1Plugin_logic_bus_rsp_payload_data;
  wire                FetchL1Plugin_logic_bus_rsp_payload_error;
  reg                 FetchL1Plugin_logic_trapPort_valid;
  reg                 FetchL1Plugin_logic_trapPort_payload_exception;
  wire       [31:0]   FetchL1Plugin_logic_trapPort_payload_tval;
  wire       [0:0]    decode_logic_trapPending;
  wire       [0:0]    DispatchPlugin_logic_trapPendings;
  wire       [0:0]    execute_lane0_logic_trapPending;
  wire                early0_IntAluPlugin_logic_wb_valid;
  wire       [31:0]   early0_IntAluPlugin_logic_wb_payload;
  (* keep , syn_keep *) reg        [31:0]   early0_IntAluPlugin_logic_alu_bitwise /* synthesis syn_keep = 1 */ ;
  wire       [31:0]   early0_IntAluPlugin_logic_alu_result;
  wire                early0_BarrelShifterPlugin_logic_wb_valid;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_wb_payload;
  wire       [4:0]    early0_BarrelShifterPlugin_logic_shift_amplitude;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_shift_reversed;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_shift_shifted;
  wire       [31:0]   early0_BarrelShifterPlugin_logic_shift_patched;
  wire                early0_BranchPlugin_logic_wb_valid;
  wire       [31:0]   early0_BranchPlugin_logic_wb_payload;
  wire                early0_BranchPlugin_logic_pcPort_valid;
  wire                early0_BranchPlugin_logic_pcPort_payload_fault;
  wire       [31:0]   early0_BranchPlugin_logic_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid;
  wire                early0_BranchPlugin_logic_historyPort_valid;
  wire       [11:0]   early0_BranchPlugin_logic_historyPort_payload_history;
  wire                early0_BranchPlugin_logic_flushPort_valid;
  wire                CfuPlugin_logic_wb_valid;
  wire       [31:0]   CfuPlugin_logic_wb_payload;
  reg                 CfuPlugin_logic_en;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3;
  reg        [2:0]    CfuPlugin_logic_csr_stateId;
  reg        [3:0]    CfuPlugin_logic_csr_cfuIndex;
  wire                CfuPlugin_logic_onFork_schedule;
  wire                CfuPlugin_logic_onFork_hold;
  reg                 CfuPlugin_logic_onFork_fired;
  wire                CfuPlugin_logic_bus_cmd_fire;
  wire                when_CfuPlugin_l147;
  wire                CfuPlugin_logic_onFork_freezeIt;
  reg                 LsuPlugin_logic_events_waiting;
  reg                 LsuPlugin_logic_trapPort_valid;
  reg                 LsuPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   LsuPlugin_logic_trapPort_payload_tval;
  wire                LsuL1_lockPort_valid;
  wire       [31:0]   LsuL1_lockPort_address;
  reg                 LsuL1_ackUnlock;
  wire                LsuL1Plugin_logic_events_loadAccess;
  wire                LsuL1Plugin_logic_events_loadMiss;
  wire                early0_MulPlugin_logic_formatBus_valid;
  wire       [31:0]   early0_MulPlugin_logic_formatBus_payload;
  wire                execute_lane0_ctrls_3_upIsCancel;
  wire                execute_lane0_ctrls_3_downIsCancel;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1;
  reg        [60:0]   _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1;
  reg        [2:0]    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2;
  wire                execute_lane0_ctrls_4_upIsCancel;
  wire                execute_lane0_ctrls_4_downIsCancel;
  reg        [65:0]   _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0;
  reg        [65:0]   _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1;
  wire                early0_DivPlugin_logic_formatBus_valid;
  wire       [31:0]   early0_DivPlugin_logic_formatBus_payload;
  reg                 early0_DivPlugin_logic_processing_divRevertResult;
  reg                 early0_DivPlugin_logic_processing_cmdSent;
  wire                early0_DivPlugin_logic_processing_div_io_cmd_fire;
  wire                early0_DivPlugin_logic_processing_request;
  wire       [31:0]   early0_DivPlugin_logic_processing_a;
  wire       [31:0]   early0_DivPlugin_logic_processing_b;
  reg                 early0_DivPlugin_logic_processing_unscheduleRequest;
  wire                early0_DivPlugin_logic_processing_freeze;
  wire       [31:0]   early0_DivPlugin_logic_processing_selected;
  wire       [31:0]   _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
  wire                CsrAccessPlugin_logic_wbWi_valid;
  wire       [31:0]   CsrAccessPlugin_logic_wbWi_payload;
  reg                 CsrAccessPlugin_logic_flushPort_valid;
  reg                 TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid;
  reg                 TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready;
  reg                 TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid;
  wire                TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready;
  reg                 early0_EnvPlugin_logic_trapPort_valid;
  reg                 early0_EnvPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   early0_EnvPlugin_logic_trapPort_payload_tval;
  reg        [3:0]    early0_EnvPlugin_logic_trapPort_payload_code;
  reg        [2:0]    early0_EnvPlugin_logic_trapPort_payload_arg;
  reg                 early0_EnvPlugin_logic_flushPort_valid;
  wire                WhiteboxerPlugin_logic_fetch_fire;
  wire       [31:0]   PrivilegedPlugin_api_lsuTriggerBus_virtual;
  wire       [1:0]    PrivilegedPlugin_api_lsuTriggerBus_size;
  wire                PrivilegedPlugin_api_harts_0_allowInterrupts;
  wire                PrivilegedPlugin_api_harts_0_allowException;
  wire                PrivilegedPlugin_api_harts_0_allowEbreakException;
  wire                PrivilegedPlugin_api_harts_0_fpuEnable;
  reg        [3:0]    CsrAccessPlugin_bus_decode_trapCode;
  wire                CsrAccessPlugin_bus_read_valid;
  wire                CsrAccessPlugin_bus_read_moving;
  wire       [11:0]   CsrAccessPlugin_bus_read_address;
  reg                 CsrAccessPlugin_bus_read_halt;
  reg        [31:0]   CsrAccessPlugin_bus_read_toWriteBits;
  wire       [31:0]   CsrAccessPlugin_bus_read_data;
  wire                CsrAccessPlugin_bus_write_valid;
  wire                CsrAccessPlugin_bus_write_moving;
  reg                 CsrAccessPlugin_bus_write_halt;
  reg        [31:0]   CsrAccessPlugin_bus_write_bits;
  wire       [11:0]   CsrAccessPlugin_bus_write_address;
  reg        [3:0]    FetchL1Plugin_logic_trapPort_payload_code;
  reg        [2:0]    FetchL1Plugin_logic_trapPort_payload_arg;
  wire                FetchL1Plugin_logic_events_access;
  wire                FetchL1Plugin_logic_events_miss;
  wire                FetchL1Plugin_logic_events_waiting;
  wire                FetchL1Plugin_logic_banks_0_write_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_0_write_payload_address;
  wire       [63:0]   FetchL1Plugin_logic_banks_0_write_payload_data;
  wire                FetchL1Plugin_logic_banks_0_read_cmd_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchL1Plugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_banks_1_write_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_1_write_payload_address;
  wire       [63:0]   FetchL1Plugin_logic_banks_1_write_payload_data;
  wire                FetchL1Plugin_logic_banks_1_read_cmd_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchL1Plugin_logic_banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_banks_2_write_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_2_write_payload_address;
  wire       [63:0]   FetchL1Plugin_logic_banks_2_write_payload_data;
  wire                FetchL1Plugin_logic_banks_2_read_cmd_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_2_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchL1Plugin_logic_banks_2_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_banks_3_write_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_3_write_payload_address;
  wire       [63:0]   FetchL1Plugin_logic_banks_3_write_payload_data;
  wire                FetchL1Plugin_logic_banks_3_read_cmd_valid;
  wire       [8:0]    FetchL1Plugin_logic_banks_3_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   FetchL1Plugin_logic_banks_3_read_rsp /* synthesis syn_keep = 1 */ ;
  reg        [3:0]    FetchL1Plugin_logic_waysWrite_mask;
  reg        [5:0]    FetchL1Plugin_logic_waysWrite_address;
  reg                 FetchL1Plugin_logic_waysWrite_tag_loaded;
  reg                 FetchL1Plugin_logic_waysWrite_tag_error;
  reg        [19:0]   FetchL1Plugin_logic_waysWrite_tag_address;
  wire                FetchL1Plugin_logic_ways_0_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_0_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_0_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_0_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_0_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded;
  wire                FetchL1Plugin_logic_ways_1_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_1_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_1_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_1_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_1_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded;
  wire                FetchL1Plugin_logic_ways_2_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_2_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_2_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_2_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_2_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_2_read_rsp_loaded;
  wire                FetchL1Plugin_logic_ways_3_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_ways_3_read_cmd_payload;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_3_read_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                FetchL1Plugin_logic_ways_3_read_rsp_error /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   FetchL1Plugin_logic_ways_3_read_rsp_address /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_FetchL1Plugin_logic_ways_3_read_rsp_loaded;
  reg                 FetchL1Plugin_logic_plru_write_valid;
  reg        [5:0]    FetchL1Plugin_logic_plru_write_payload_address;
  reg        [0:0]    FetchL1Plugin_logic_plru_write_payload_data_0;
  reg        [1:0]    FetchL1Plugin_logic_plru_write_payload_data_1;
  wire                FetchL1Plugin_logic_plru_read_cmd_valid;
  wire       [5:0]    FetchL1Plugin_logic_plru_read_cmd_payload;
  (* keep , syn_keep *) wire       [0:0]    FetchL1Plugin_logic_plru_read_rsp_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [1:0]    FetchL1Plugin_logic_plru_read_rsp_1 /* synthesis syn_keep = 1 */ ;
  wire       [2:0]    _zz_FetchL1Plugin_logic_plru_read_rsp_0;
  wire                FetchL1Plugin_logic_invalidate_cmd_valid;
  wire                FetchL1Plugin_logic_invalidate_cmd_ready;
  reg                 FetchL1Plugin_logic_invalidate_canStart;
  reg        [6:0]    FetchL1Plugin_logic_invalidate_counter;
  wire       [6:0]    FetchL1Plugin_logic_invalidate_counterIncr;
  wire                FetchL1Plugin_logic_invalidate_done;
  wire                FetchL1Plugin_logic_invalidate_last;
  reg                 FetchL1Plugin_logic_invalidate_firstEver;
  wire                when_FetchL1Plugin_l204;
  wire                when_FetchL1Plugin_l211;
  wire                when_FetchL1Plugin_l216;
  wire                fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217;
  reg                 FetchL1Plugin_logic_refill_start_valid;
  wire       [31:0]   FetchL1Plugin_logic_refill_start_address;
  wire       [1:0]    FetchL1Plugin_logic_refill_start_wayToAllocate;
  wire                FetchL1Plugin_logic_refill_start_isIo;
  reg                 FetchL1Plugin_logic_refill_slots_0_valid;
  reg                 FetchL1Plugin_logic_refill_slots_0_cmdSent;
  (* keep , syn_keep *) reg        [31:0]   FetchL1Plugin_logic_refill_slots_0_address /* synthesis syn_keep = 1 */ ;
  reg                 FetchL1Plugin_logic_refill_slots_0_isIo;
  reg        [1:0]    FetchL1Plugin_logic_refill_slots_0_wayToAllocate;
  reg        [0:0]    FetchL1Plugin_logic_refill_slots_0_priority;
  wire                FetchL1Plugin_logic_refill_slots_0_askCmd;
  reg        [31:0]   FetchL1Plugin_logic_refill_pushCounter;
  wire                FetchL1Plugin_logic_refill_hazard;
  wire                when_FetchL1Plugin_l255;
  wire                when_FetchL1Plugin_l268;
  wire       [0:0]    FetchL1Plugin_logic_refill_onCmd_propoedOh;
  reg                 FetchL1Plugin_logic_refill_onCmd_locked;
  wire                when_FetchL1Plugin_l276;
  reg        [0:0]    FetchL1Plugin_logic_refill_onCmd_lockedOh;
  wire       [0:0]    FetchL1Plugin_logic_refill_onCmd_oh;
  (* keep , syn_keep *) reg        [2:0]    FetchL1Plugin_logic_refill_onRsp_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                FetchL1Plugin_logic_refill_onRsp_holdHarts;
  wire                fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l297;
  reg                 FetchL1Plugin_logic_refill_onRsp_firstCycle;
  wire                FetchL1Plugin_logic_bus_rsp_fire;
  wire       [1:0]    FetchL1Plugin_logic_refill_onRsp_wayToAllocate;
  wire       [31:0]   FetchL1Plugin_logic_refill_onRsp_address;
  wire                when_FetchL1Plugin_l304;
  wire                when_FetchL1Plugin_l330;
  wire                FetchL1Plugin_logic_cmd_doIt;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_0;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_1;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_2;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_translatedHits;
  wire                FetchL1Plugin_logic_hits_w_0_indirect_bypassHits;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_0;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_1;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_2;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_translatedHits;
  wire                FetchL1Plugin_logic_hits_w_1_indirect_bypassHits;
  wire                FetchL1Plugin_logic_hits_w_2_indirect_wayTlbHits_0;
  wire                FetchL1Plugin_logic_hits_w_2_indirect_wayTlbHits_1;
  wire                FetchL1Plugin_logic_hits_w_2_indirect_wayTlbHits_2;
  wire                FetchL1Plugin_logic_hits_w_2_indirect_translatedHits;
  wire                FetchL1Plugin_logic_hits_w_2_indirect_bypassHits;
  wire                FetchL1Plugin_logic_hits_w_3_indirect_wayTlbHits_0;
  wire                FetchL1Plugin_logic_hits_w_3_indirect_wayTlbHits_1;
  wire                FetchL1Plugin_logic_hits_w_3_indirect_wayTlbHits_2;
  wire                FetchL1Plugin_logic_hits_w_3_indirect_translatedHits;
  wire                FetchL1Plugin_logic_hits_w_3_indirect_bypassHits;
  wire       [31:0]   FetchL1Plugin_logic_ctrl_pmaPort_cmd_address;
  wire                FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault;
  wire                FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0;
  wire       [1:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_1;
  wire       [1:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id;
  wire       [1:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0;
  reg        [1:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_1;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_1;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_1_stateSel;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_1_state;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_core_update_logic_1_sel;
  wire                _zz_FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id;
  wire                _zz_FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id_1;
  wire                FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid;
  wire       [5:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address;
  wire       [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0;
  wire       [1:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_1;
  reg                 FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid;
  reg        [5:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address;
  reg        [0:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0;
  reg        [1:0]    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_1;
  wire                FetchL1Plugin_logic_ctrl_dataAccessFault;
  reg                 FetchL1Plugin_logic_ctrl_trapSent;
  reg                 FetchL1Plugin_logic_ctrl_allowRefill;
  wire                when_FetchL1Plugin_l474;
  wire                when_FetchL1Plugin_l480;
  wire                when_FetchL1Plugin_l487;
  wire                when_FetchL1Plugin_l520;
  wire                when_FetchL1Plugin_l533;
  wire                when_FetchL1Plugin_l537;
  reg                 FetchL1Plugin_logic_ctrl_firstCycle;
  wire                when_FetchL1Plugin_l541;
  reg                 FetchL1Plugin_logic_ctrl_onEvents_waiting;
  wire                when_FetchL1Plugin_l549;
  wire                when_FetchL1Plugin_l558;
  wire       [2:0]    _zz_FetchL1Plugin_logic_plru_write_payload_data_0;
  reg        [3:0]    LsuPlugin_logic_trapPort_payload_code;
  reg        [2:0]    LsuPlugin_logic_trapPort_payload_arg;
  reg                 LsuPlugin_logic_flushPort_valid;
  wire       [15:0]   LsuPlugin_logic_flushPort_payload_uopId;
  wire                LsuPlugin_logic_flushPort_payload_self;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_0;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_1;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_2;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_3;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_4;
  wire                LsuPlugin_logic_frontend_defaultsDecodings_5;
  wire                LsuPlugin_logic_commitProbe_valid;
  wire       [31:0]   LsuPlugin_logic_commitProbe_payload_pc;
  wire       [31:0]   LsuPlugin_logic_commitProbe_payload_address;
  wire                LsuPlugin_logic_commitProbe_payload_load;
  wire                LsuPlugin_logic_commitProbe_payload_store;
  wire                LsuPlugin_logic_commitProbe_payload_trap;
  wire                LsuPlugin_logic_commitProbe_payload_io;
  wire                LsuPlugin_logic_commitProbe_payload_prefetchFailed;
  wire                LsuPlugin_logic_commitProbe_payload_miss;
  wire                LsuPlugin_logic_iwb_valid;
  reg        [31:0]   LsuPlugin_logic_iwb_payload;
  wire                execute_lane0_ctrls_0_upIsCancel;
  wire                execute_lane0_ctrls_0_downIsCancel;
  reg                 PrivilegedPlugin_logic_harts_0_xretAwayFromMachine;
  wire       [0:0]    PrivilegedPlugin_logic_harts_0_commitMask;
  reg                 PrivilegedPlugin_logic_harts_0_int_pending;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_privilege;
  wire                PrivilegedPlugin_logic_harts_0_withMachinePrivilege;
  wire                PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege;
  wire                PrivilegedPlugin_logic_harts_0_hartRunning;
  wire                PrivilegedPlugin_logic_harts_0_debugMode;
  wire                when_CsrService_l198;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mie;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mpie;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_m_status_mpp;
  reg        [1:0]    PrivilegedPlugin_logic_harts_0_m_status_fs;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_sd;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_tsr;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_tvm;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_tw;
  reg                 PrivilegedPlugin_logic_harts_0_m_status_mprv;
  wire                when_PrivilegedPlugin_l542;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4;
  wire                when_CsrService_l176;
  reg                 PrivilegedPlugin_logic_harts_0_m_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_harts_0_m_cause_code;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_meip;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_mtip;
  reg                 PrivilegedPlugin_logic_harts_0_m_ip_msip;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_meie;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_mtie;
  reg                 PrivilegedPlugin_logic_harts_0_m_ie_msie;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_iam;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_bp;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_eu;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_es;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_ipf;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_lpf;
  reg                 PrivilegedPlugin_logic_harts_0_m_edeleg_spf;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10;
  reg                 PrivilegedPlugin_logic_harts_0_m_ideleg_st;
  reg                 PrivilegedPlugin_logic_harts_0_m_ideleg_se;
  reg                 PrivilegedPlugin_logic_harts_0_m_ideleg_ss;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12;
  wire                _zz_when_TrapPlugin_l207;
  wire                _zz_when_TrapPlugin_l207_1;
  wire                _zz_when_TrapPlugin_l207_2;
  reg                 PrivilegedPlugin_logic_harts_0_s_cause_interrupt;
  reg        [3:0]    PrivilegedPlugin_logic_harts_0_s_cause_code;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13;
  reg                 PrivilegedPlugin_logic_harts_0_s_status_sie;
  reg                 PrivilegedPlugin_logic_harts_0_s_status_spie;
  reg        [0:0]    PrivilegedPlugin_logic_harts_0_s_status_spp;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_seipSoft;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_seipInput;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_seipOr;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_stip;
  reg                 PrivilegedPlugin_logic_harts_0_s_ip_ssip;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_seipMasked;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_stipMasked;
  wire                PrivilegedPlugin_logic_harts_0_s_ip_ssipMasked;
  reg                 PrivilegedPlugin_logic_harts_0_s_ie_seie;
  reg                 PrivilegedPlugin_logic_harts_0_s_ie_stie;
  reg                 PrivilegedPlugin_logic_harts_0_s_ie_ssie;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16;
  wire                _zz_when_TrapPlugin_l207_3;
  wire                _zz_when_TrapPlugin_l207_4;
  wire                _zz_when_TrapPlugin_l207_5;
  wire       [1:0]    PrivilegedPlugin_logic_defaultTrap_csrPrivilege;
  wire                PrivilegedPlugin_logic_defaultTrap_csrReadOnly;
  wire                when_PrivilegedPlugin_l689;
  wire                GSharePlugin_logic_mem_write_valid;
  wire       [13:0]   GSharePlugin_logic_mem_write_payload_address;
  wire       [1:0]    GSharePlugin_logic_mem_write_payload_data_0;
  wire       [13:0]   _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
  wire                when_GSharePlugin_l88;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_push;
  reg        [1:0]    BtbPlugin_logic_ras_ptr_pop;
  reg                 BtbPlugin_logic_ras_ptr_pushIt;
  reg                 BtbPlugin_logic_ras_ptr_popIt;
  wire                BtbPlugin_logic_ras_readIt;
  reg        [29:0]   BtbPlugin_logic_ras_read;
  wire                BtbPlugin_logic_ras_write_valid;
  wire       [1:0]    BtbPlugin_logic_ras_write_payload_address;
  reg        [29:0]   BtbPlugin_logic_ras_write_payload_data;
  reg                 BtbPlugin_logic_memWrite_valid;
  reg        [8:0]    BtbPlugin_logic_memWrite_payload_address;
  reg        [15:0]   BtbPlugin_logic_memWrite_payload_data_0_hash;
  wire       [29:0]   BtbPlugin_logic_memWrite_payload_data_0_pcTarget;
  reg                 BtbPlugin_logic_memWrite_payload_data_0_isBranch;
  reg                 BtbPlugin_logic_memWrite_payload_data_0_isPush;
  reg                 BtbPlugin_logic_memWrite_payload_data_0_isPop;
  reg        [0:0]    BtbPlugin_logic_memWrite_payload_mask;
  wire                BtbPlugin_logic_memRead_cmd_valid;
  wire       [8:0]    BtbPlugin_logic_memRead_cmd_payload;
  wire       [15:0]   BtbPlugin_logic_memRead_rsp_0_hash;
  wire       [29:0]   BtbPlugin_logic_memRead_rsp_0_pcTarget;
  wire                BtbPlugin_logic_memRead_rsp_0_isBranch;
  wire                BtbPlugin_logic_memRead_rsp_0_isPush;
  wire                BtbPlugin_logic_memRead_rsp_0_isPop;
  wire                BtbPlugin_logic_memDp_wp_valid;
  wire       [8:0]    BtbPlugin_logic_memDp_wp_payload_address;
  wire       [15:0]   BtbPlugin_logic_memDp_wp_payload_data_0_hash;
  wire       [29:0]   BtbPlugin_logic_memDp_wp_payload_data_0_pcTarget;
  wire                BtbPlugin_logic_memDp_wp_payload_data_0_isBranch;
  wire                BtbPlugin_logic_memDp_wp_payload_data_0_isPush;
  wire                BtbPlugin_logic_memDp_wp_payload_data_0_isPop;
  wire       [0:0]    BtbPlugin_logic_memDp_wp_payload_mask;
  wire                BtbPlugin_logic_memDp_rp_cmd_valid;
  wire       [8:0]    BtbPlugin_logic_memDp_rp_cmd_payload;
  wire       [15:0]   BtbPlugin_logic_memDp_rp_rsp_0_hash;
  wire       [29:0]   BtbPlugin_logic_memDp_rp_rsp_0_pcTarget;
  wire                BtbPlugin_logic_memDp_rp_rsp_0_isBranch;
  wire                BtbPlugin_logic_memDp_rp_rsp_0_isPush;
  wire                BtbPlugin_logic_memDp_rp_rsp_0_isPop;
  wire       [48:0]   _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash;
  wire       [9:0]    WhiteboxerPlugin_logic_fetch_fetchId;
  wire                WhiteboxerPlugin_logic_decodes_0_fire;
  reg                 decode_ctrls_0_up_LANE_SEL_0_regNext;
  wire                when_CtrlLaneApi_l50;
  wire                WhiteboxerPlugin_logic_decodes_0_spawn;
  wire       [63:0]   WhiteboxerPlugin_logic_decodes_0_pc;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_0_fetchId;
  wire       [9:0]    WhiteboxerPlugin_logic_decodes_0_decodeId;
  wire       [15:0]   early0_BranchPlugin_logic_flushPort_payload_uopId;
  wire                early0_BranchPlugin_logic_flushPort_payload_self;
  reg                 early0_BranchPlugin_logic_trapPort_valid;
  wire                early0_BranchPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   early0_BranchPlugin_logic_trapPort_payload_tval;
  wire       [3:0]    early0_BranchPlugin_logic_trapPort_payload_code;
  wire       [2:0]    early0_BranchPlugin_logic_trapPort_payload_arg;
  wire       [15:0]   CsrAccessPlugin_logic_flushPort_payload_uopId;
  wire                CsrAccessPlugin_logic_flushPort_payload_self;
  reg                 CsrAccessPlugin_logic_trapPort_valid;
  reg                 CsrAccessPlugin_logic_trapPort_payload_exception;
  wire       [31:0]   CsrAccessPlugin_logic_trapPort_payload_tval;
  reg        [3:0]    CsrAccessPlugin_logic_trapPort_payload_code;
  wire       [2:0]    CsrAccessPlugin_logic_trapPort_payload_arg;
  wire       [15:0]   early0_EnvPlugin_logic_flushPort_payload_uopId;
  wire                early0_EnvPlugin_logic_flushPort_payload_self;
  wire       [1:0]    early0_EnvPlugin_logic_exe_privilege;
  wire       [0:0]    MmuPlugin_logic_satpModeWrite;
  reg                 DecoderPlugin_logic_forgetPort_valid;
  reg        [31:0]   DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice;
  wire       [0:0]    PerformanceCounterPlugin_logic_commitMask;
  reg                 PerformanceCounterPlugin_logic_ignoreNextCommit;
  wire                when_PerformanceCounterPlugin_l45;
  wire       [0:0]    PerformanceCounterPlugin_logic_commitCount;
  wire                PerformanceCounterPlugin_logic_eventCycles;
  wire                PerformanceCounterPlugin_logic_eventInstructions_0;
  reg        [7:0]    PerformanceCounterPlugin_logic_counters_cycle_value;
  wire                PerformanceCounterPlugin_logic_counters_cycle_needFlush;
  reg                 PerformanceCounterPlugin_logic_counters_cycle_mcounteren;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17;
  reg                 PerformanceCounterPlugin_logic_counters_cycle_scounteren;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18;
  reg                 PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit;
  wire                _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19;
  reg        [7:0]    PerformanceCounterPlugin_logic_counters_instret_value;
  wire                PerformanceCounterPlugin_logic_counters_instret_needFlush;
  reg                 PerformanceCounterPlugin_logic_counters_instret_mcounteren;
  reg                 PerformanceCounterPlugin_logic_counters_instret_scounteren;
  reg                 PerformanceCounterPlugin_logic_counters_instret_mcountinhibit;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_counters_instret_value;
  wire                execute_lane0_ctrls_1_upIsCancel;
  wire                execute_lane0_ctrls_1_downIsCancel;
  reg        [31:0]   _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  reg        [31:0]   _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  reg        [31:0]   early0_SrcPlugin_logic_addsub_combined_rs2Patched;
  wire                lane0_IntFormatPlugin_logic_stages_0_wb_valid;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_0_wb_payload;
  wire       [1:0]    lane0_IntFormatPlugin_logic_stages_0_hits;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_0_raw;
  wire                lane0_IntFormatPlugin_logic_stages_1_wb_valid;
  reg        [31:0]   lane0_IntFormatPlugin_logic_stages_1_wb_payload;
  wire       [1:0]    lane0_IntFormatPlugin_logic_stages_1_hits;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_1_raw;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_sels_0;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_0_doIt;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_0;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_1;
  reg                 _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value;
  wire                lane0_IntFormatPlugin_logic_stages_1_segments_1_doIt;
  wire                lane0_IntFormatPlugin_logic_stages_2_wb_valid;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_2_wb_payload;
  wire       [1:0]    lane0_IntFormatPlugin_logic_stages_2_hits;
  wire       [31:0]   lane0_IntFormatPlugin_logic_stages_2_raw;
  reg        [31:0]   early0_BranchPlugin_pcCalc_target_a;
  reg        [31:0]   early0_BranchPlugin_pcCalc_target_b;
  wire       [1:0]    early0_BranchPlugin_pcCalc_slices;
  wire       [0:0]    AlignerPlugin_logic_maskGen_frontMasks_0;
  wire       [0:0]    AlignerPlugin_logic_maskGen_backMasks_0;
  wire       [31:0]   AlignerPlugin_logic_slices_data_0;
  wire       [0:0]    AlignerPlugin_logic_slices_mask;
  wire       [0:0]    AlignerPlugin_logic_slices_last;
  wire       [31:0]   AlignerPlugin_logic_slicesInstructions_0;
  reg        [0:0]    AlignerPlugin_logic_scanners_0_usageMask;
  wire                AlignerPlugin_logic_scanners_0_checker_0_required;
  wire                AlignerPlugin_logic_scanners_0_checker_0_last;
  wire                AlignerPlugin_logic_scanners_0_checker_0_redo;
  wire                AlignerPlugin_logic_scanners_0_checker_0_present;
  wire                AlignerPlugin_logic_scanners_0_checker_0_valid;
  wire                AlignerPlugin_logic_scanners_0_redo;
  wire                AlignerPlugin_logic_scanners_0_valid;
  wire       [0:0]    AlignerPlugin_logic_usedMask_0;
  wire       [0:0]    AlignerPlugin_logic_usedMask_1;
  wire                AlignerPlugin_logic_extractors_0_first;
  wire       [0:0]    AlignerPlugin_logic_extractors_0_usableMask;
  wire                AlignerPlugin_logic_extractors_0_usableMask_bools_0;
  wire       [0:0]    _zz_AlignerPlugin_logic_extractors_0_slicesOh;
  wire       [0:0]    AlignerPlugin_logic_extractors_0_slicesOh;
  reg                 AlignerPlugin_logic_extractors_0_redo;
  wire       [0:0]    AlignerPlugin_logic_extractors_0_localMask;
  reg        [0:0]    AlignerPlugin_logic_extractors_0_usageMask;
  reg                 AlignerPlugin_logic_extractors_0_valid;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_ctx_pc;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_ctx_instruction;
  wire       [9:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID;
  wire       [1:0]    AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [11:0]   AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY;
  wire       [0:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  wire       [0:0]    AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  wire       [31:0]   AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC;
  wire                AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED;
  wire                AlignerPlugin_logic_extractors_0_ctx_trap;
  wire                when_AlignerPlugin_l160;
  reg        [9:0]    AlignerPlugin_logic_feeder_harts_0_dopId;
  wire                when_AlignerPlugin_l171;
  wire                AlignerPlugin_logic_feeder_lanes_0_valid;
  wire                AlignerPlugin_logic_feeder_lanes_0_isRvc;
  wire                AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction;
  reg        [0:0]    AlignerPlugin_logic_nobuffer_mask;
  wire       [0:0]    AlignerPlugin_logic_nobuffer_remaningMask;
  wire                when_AlignerPlugin_l292;
  wire       [2:0]    CfuPlugin_logic_onFork_functionsIds_0;
  wire       [2:0]    CfuPlugin_logic_onFork_functionsIds_1;
  reg        [31:0]   _zz_CfuPlugin_logic_bus_cmd_payload_inputs_1;
  wire                CfuPlugin_logic_bus_rsp_toFlow_valid;
  wire       [31:0]   CfuPlugin_logic_bus_rsp_toFlow_payload_outputs_0;
  wire                CfuPlugin_logic_onJoin_busRspStream_valid;
  wire                CfuPlugin_logic_onJoin_busRspStream_ready;
  wire       [31:0]   CfuPlugin_logic_onJoin_busRspStream_payload_outputs_0;
  wire                CfuPlugin_logic_onJoin_freezeIt;
  wire                LsuPlugin_logic_bus_cmd_valid;
  wire                LsuPlugin_logic_bus_cmd_ready;
  wire                LsuPlugin_logic_bus_cmd_payload_write;
  wire       [31:0]   LsuPlugin_logic_bus_cmd_payload_address;
  wire       [31:0]   LsuPlugin_logic_bus_cmd_payload_data;
  wire       [1:0]    LsuPlugin_logic_bus_cmd_payload_size;
  wire       [3:0]    LsuPlugin_logic_bus_cmd_payload_mask;
  wire                LsuPlugin_logic_bus_cmd_payload_io;
  wire                LsuPlugin_logic_bus_cmd_payload_fromHart;
  wire       [15:0]   LsuPlugin_logic_bus_cmd_payload_uopId;
  wire                LsuPlugin_logic_bus_rsp_valid;
  wire                LsuPlugin_logic_bus_rsp_payload_error;
  wire       [31:0]   LsuPlugin_logic_bus_rsp_payload_data;
  wire                LsuPlugin_logic_flusher_wantExit;
  reg                 LsuPlugin_logic_flusher_wantStart;
  wire                LsuPlugin_logic_flusher_wantKill;
  reg        [6:0]    LsuPlugin_logic_flusher_cmdCounter;
  wire                LsuPlugin_logic_flusher_inflight;
  wire       [1:0]    early0_EnvPlugin_logic_exe_xretPriv;
  reg                 early0_EnvPlugin_logic_exe_commit;
  wire                early0_EnvPlugin_logic_exe_retKo;
  wire                early0_EnvPlugin_logic_exe_vmaKo;
  wire                when_EnvPlugin_l86;
  wire                when_EnvPlugin_l95;
  wire                when_EnvPlugin_l110;
  wire                when_EnvPlugin_l119;
  wire                when_EnvPlugin_l123;
  reg                 PerformanceCounterPlugin_logic_readPort_valid;
  wire                PerformanceCounterPlugin_logic_readPort_ready;
  wire       [3:0]    PerformanceCounterPlugin_logic_readPort_address;
  wire       [31:0]   PerformanceCounterPlugin_logic_readPort_data;
  reg                 PerformanceCounterPlugin_logic_writePort_valid;
  wire                PerformanceCounterPlugin_logic_writePort_ready;
  wire       [3:0]    PerformanceCounterPlugin_logic_writePort_address;
  reg        [31:0]   PerformanceCounterPlugin_logic_writePort_data;
  wire                CsrRamPlugin_setup_initPort_valid;
  wire                CsrRamPlugin_setup_initPort_ready;
  wire       [3:0]    CsrRamPlugin_setup_initPort_address;
  wire       [31:0]   CsrRamPlugin_setup_initPort_data;
  wire                early0_BranchPlugin_logic_alu_expectedMsb;
  wire       [2:0]    switch_Misc_l242;
  reg                 _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  reg                 _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  wire                early0_BranchPlugin_logic_jumpLogic_wrongCond;
  wire                early0_BranchPlugin_logic_jumpLogic_needFix;
  wire                early0_BranchPlugin_logic_jumpLogic_doIt;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_fetched;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_next;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_history_shifter;
  wire                when_BranchPlugin_l218;
  wire                when_BranchPlugin_l251;
  wire                early0_BranchPlugin_logic_jumpLogic_rdLink;
  wire                early0_BranchPlugin_logic_jumpLogic_rs1Link;
  wire                early0_BranchPlugin_logic_jumpLogic_rdEquRs1;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_valid;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_ready;
  wire       [31:0]   early0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  wire       [31:0]   early0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  wire       [15:0]   early0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  wire       [1:0]    early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire                CsrRamPlugin_csrMapper_read_valid;
  wire                CsrRamPlugin_csrMapper_read_ready;
  wire       [3:0]    CsrRamPlugin_csrMapper_read_address;
  wire       [31:0]   CsrRamPlugin_csrMapper_read_data;
  wire                CsrRamPlugin_csrMapper_write_valid;
  wire                CsrRamPlugin_csrMapper_write_ready;
  wire       [3:0]    CsrRamPlugin_csrMapper_write_address;
  wire       [31:0]   CsrRamPlugin_csrMapper_write_data;
  wire                LearnPlugin_logic_learn_valid;
  wire       [31:0]   LearnPlugin_logic_learn_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_learn_payload_pcTarget;
  wire                LearnPlugin_logic_learn_payload_taken;
  wire                LearnPlugin_logic_learn_payload_isBranch;
  wire                LearnPlugin_logic_learn_payload_isPush;
  wire                LearnPlugin_logic_learn_payload_isPop;
  wire                LearnPlugin_logic_learn_payload_wasWrong;
  wire                LearnPlugin_logic_learn_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_learn_payload_history;
  wire       [15:0]   LearnPlugin_logic_learn_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire                LearnPlugin_logic_buffered_0_valid;
  wire                LearnPlugin_logic_buffered_0_ready;
  wire       [31:0]   LearnPlugin_logic_buffered_0_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_buffered_0_payload_pcTarget;
  wire                LearnPlugin_logic_buffered_0_payload_taken;
  wire                LearnPlugin_logic_buffered_0_payload_isBranch;
  wire                LearnPlugin_logic_buffered_0_payload_isPush;
  wire                LearnPlugin_logic_buffered_0_payload_isPop;
  wire                LearnPlugin_logic_buffered_0_payload_wasWrong;
  wire                LearnPlugin_logic_buffered_0_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_buffered_0_payload_history;
  wire       [15:0]   LearnPlugin_logic_buffered_0_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire                LearnPlugin_logic_arbitrated_valid;
  wire                LearnPlugin_logic_arbitrated_ready;
  wire       [31:0]   LearnPlugin_logic_arbitrated_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_arbitrated_payload_pcTarget;
  wire                LearnPlugin_logic_arbitrated_payload_taken;
  wire                LearnPlugin_logic_arbitrated_payload_isBranch;
  wire                LearnPlugin_logic_arbitrated_payload_isPush;
  wire                LearnPlugin_logic_arbitrated_payload_isPop;
  wire                LearnPlugin_logic_arbitrated_payload_wasWrong;
  wire                LearnPlugin_logic_arbitrated_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_arbitrated_payload_history;
  wire       [15:0]   LearnPlugin_logic_arbitrated_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire                LearnPlugin_logic_arbitrated_toFlow_valid;
  wire       [31:0]   LearnPlugin_logic_arbitrated_toFlow_payload_pcOnLastSlice;
  wire       [31:0]   LearnPlugin_logic_arbitrated_toFlow_payload_pcTarget;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_taken;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_isBranch;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_isPush;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_isPop;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_wasWrong;
  wire                LearnPlugin_logic_arbitrated_toFlow_payload_badPredictedTarget;
  wire       [11:0]   LearnPlugin_logic_arbitrated_toFlow_payload_history;
  wire       [15:0]   LearnPlugin_logic_arbitrated_toFlow_payload_uopId;
  wire       [1:0]    LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  reg        [15:0]   DecoderPlugin_logic_harts_0_uopId;
  wire                when_DecoderPlugin_l143;
  wire       [0:0]    DecoderPlugin_logic_interrupt_async;
  wire                when_DecoderPlugin_l151;
  reg        [0:0]    DecoderPlugin_logic_interrupt_buffered;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  wire                _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  wire                when_CfuPlugin_l115;
  wire                DecoderPlugin_logic_laneLogic_0_interruptPending;
  reg                 DecoderPlugin_logic_laneLogic_0_trapPort_valid;
  reg                 DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception;
  wire       [31:0]   DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval;
  reg        [3:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_code;
  wire       [2:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg;
  wire       [0:0]    DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge;
  wire                DecoderPlugin_logic_laneLogic_0_fixer_isJb;
  wire                DecoderPlugin_logic_laneLogic_0_fixer_doIt;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap;
  wire                DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit;
  reg                 decode_ctrls_1_up_LANE_SEL_0_regNext;
  wire                when_CtrlLaneApi_l50_1;
  wire                when_DecoderPlugin_l229;
  wire                DecoderPlugin_logic_laneLogic_0_flushPort_valid;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId;
  wire                DecoderPlugin_logic_laneLogic_0_flushPort_payload_self;
  wire                when_DecoderPlugin_l247;
  wire       [15:0]   DecoderPlugin_logic_laneLogic_0_uopIdBase;
  wire                DispatchPlugin_logic_candidates_0_ctx_valid;
  reg        [0:0]    DispatchPlugin_logic_candidates_0_ctx_laneLayerHits;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_uop;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  wire       [1:0]    DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  wire       [11:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  wire       [31:0]   DispatchPlugin_logic_candidates_0_ctx_hm_PC;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_TRAP;
  wire       [15:0]   DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE;
  wire       [4:0]    DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  wire                DispatchPlugin_logic_candidates_0_fire;
  wire                DispatchPlugin_logic_candidates_0_cancel;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_rsHazards;
  wire       [0:0]    DispatchPlugin_logic_candidates_0_reservationHazards;
  wire                DispatchPlugin_logic_candidates_0_flushHazards;
  wire                DispatchPlugin_logic_candidates_0_fenceOlderHazards;
  wire                DispatchPlugin_logic_candidates_0_moving;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard;
  wire                DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard;
  wire                DispatchPlugin_logic_reservationChecker_0_onLl_0_hit;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0;
  wire                DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1;
  wire                DispatchPlugin_logic_flushChecker_0_oldersHazard;
  wire       [0:0]    DispatchPlugin_logic_fenceChecker_olderInflights;
  wire                DispatchPlugin_logic_feeds_0_sending;
  reg                 DispatchPlugin_logic_feeds_0_sent;
  wire                when_DispatchPlugin_l368;
  wire       [0:0]    DispatchPlugin_logic_scheduler_eusFree_0;
  wire       [0:0]    DispatchPlugin_logic_scheduler_eusFree_1;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_0;
  wire       [0:0]    DispatchPlugin_logic_scheduler_hartFree_1;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_candHazard;
  wire       [0:0]    DispatchPlugin_logic_scheduler_arbiters_0_layersHits;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0;
  wire       [0:0]    _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  wire       [0:0]    DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  wire       [0:0]    DispatchPlugin_logic_scheduler_arbiters_0_eusOh;
  wire                DispatchPlugin_logic_scheduler_arbiters_0_doIt;
  wire       [0:0]    DispatchPlugin_logic_inserter_0_oh;
  wire                DispatchPlugin_logic_inserter_0_trap;
  wire                when_DispatchPlugin_l439;
  wire       [0:0]    DispatchPlugin_logic_inserter_0_layerOhUnfiltred;
  wire                DispatchPlugin_logic_inserter_0_layer_0_1;
  wire                DispatchPlugin_logic_events_frontendStall;
  wire                DispatchPlugin_logic_events_backendStall;
  wire       [3:0]    CsrRamPlugin_csrMapper_ramAddress;
  wire       [11:0]   _zz_CsrRamPlugin_csrMapper_ramAddress;
  reg                 CsrRamPlugin_csrMapper_withRead;
  wire                when_CsrRamPlugin_l85;
  reg                 CsrRamPlugin_csrMapper_doWrite;
  reg                 CsrRamPlugin_csrMapper_fired;
  wire                when_CsrRamPlugin_l92;
  wire                when_CsrRamPlugin_l96;
  wire       [13:0]   _zz_GSharePlugin_logic_onLearn_hash;
  wire       [13:0]   GSharePlugin_logic_onLearn_hash;
  wire       [1:0]    GSharePlugin_logic_onLearn_updated_0;
  wire       [1:0]    GSharePlugin_logic_onLearn_incrValue;
  reg                 GSharePlugin_logic_onLearn_overflow;
  wire                when_GSharePlugin_l107;
  wire       [15:0]   BtbPlugin_logic_onLearn_hash;
  wire       [1:0]    lane0_integer_WriteBackPlugin_logic_stages_0_hits;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  wire                lane0_integer_WriteBackPlugin_logic_stages_0_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  wire       [0:0]    lane0_integer_WriteBackPlugin_logic_stages_1_hits;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_1_muxed;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_1_merged;
  wire                lane0_integer_WriteBackPlugin_logic_stages_1_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  wire       [1:0]    lane0_integer_WriteBackPlugin_logic_stages_2_hits;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_2_muxed;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_2_merged;
  wire                lane0_integer_WriteBackPlugin_logic_stages_2_write_valid;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  wire                lane0_integer_WriteBackPlugin_logic_write_port_valid;
  wire       [4:0]    lane0_integer_WriteBackPlugin_logic_write_port_address;
  wire       [31:0]   lane0_integer_WriteBackPlugin_logic_write_port_data;
  wire       [15:0]   lane0_integer_WriteBackPlugin_logic_write_port_uopId;
  wire                _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  wire                _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1;
  wire                _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2;
  wire                TrapPlugin_logic_initHold;
  reg                 decode_ctrls_1_up_LANE_SEL_0_regNext_1;
  wire                when_CtrlLaneApi_l50_2;
  wire                WhiteboxerPlugin_logic_serializeds_0_fire;
  wire       [9:0]    WhiteboxerPlugin_logic_serializeds_0_decodeId;
  wire       [15:0]   WhiteboxerPlugin_logic_serializeds_0_microOpId;
  wire       [31:0]   WhiteboxerPlugin_logic_serializeds_0_microOp;
  reg                 execute_ctrl0_down_LANE_SEL_lane0_regNext;
  wire                when_CtrlLaneApi_l50_3;
  wire                WhiteboxerPlugin_logic_dispatches_0_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_dispatches_0_microOpId;
  reg                 execute_ctrl2_down_LANE_SEL_lane0_regNext;
  wire                when_CtrlLaneApi_l50_4;
  wire                WhiteboxerPlugin_logic_executes_0_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_executes_0_microOpId;
  wire                WhiteboxerPlugin_logic_csr_access_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_csr_access_payload_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_csr_access_payload_address;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_access_payload_write;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_access_payload_read;
  wire                WhiteboxerPlugin_logic_csr_access_payload_writeDone;
  wire                WhiteboxerPlugin_logic_csr_access_payload_readDone;
  wire       [15:0]   BtbPlugin_logic_onForget_hash;
  wire                fetch_logic_ctrls_0_haltRequest_BtbPlugin_l200;
  wire       [0:0]    BtbPlugin_logic_predictions;
  wire       [0:0]    BtbPlugin_logic_applyIt_chunksMask;
  wire       [0:0]    BtbPlugin_logic_applyIt_chunksTakenOh;
  wire                BtbPlugin_logic_applyIt_needIt;
  reg                 BtbPlugin_logic_applyIt_correctionSent;
  wire                when_BtbPlugin_l233;
  wire                BtbPlugin_logic_applyIt_doIt;
  wire       [15:0]   BtbPlugin_logic_applyIt_entry_hash;
  wire       [29:0]   BtbPlugin_logic_applyIt_entry_pcTarget;
  wire                BtbPlugin_logic_applyIt_entry_isBranch;
  wire                BtbPlugin_logic_applyIt_entry_isPush;
  wire                BtbPlugin_logic_applyIt_entry_isPop;
  reg        [29:0]   BtbPlugin_logic_applyIt_pcTarget;
  wire                BtbPlugin_logic_applyIt_rasLogic_pushValid;
  wire       [31:0]   BtbPlugin_logic_applyIt_rasLogic_pushPc;
  wire                when_BtbPlugin_l246;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_0_history;
  wire                BtbPlugin_logic_applyIt_history_layers_0_valid;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layers_1_history;
  wire                BtbPlugin_logic_applyIt_history_layers_1_valid;
  wire                BtbPlugin_logic_applyIt_history_layersLogic_0_doIt;
  wire       [11:0]   BtbPlugin_logic_applyIt_history_layersLogic_0_shifted;
  reg                 TrapPlugin_logic_harts_0_crsPorts_read_valid;
  wire                TrapPlugin_logic_harts_0_crsPorts_read_ready;
  reg        [3:0]    TrapPlugin_logic_harts_0_crsPorts_read_address;
  wire       [31:0]   TrapPlugin_logic_harts_0_crsPorts_read_data;
  wire                AlignerPlugin_logic_nobuffer_flushIt;
  wire                when_AlignerPlugin_l298;
  wire                decode_logic_flushes_0_onLanes_0_doIt;
  wire                decode_logic_flushes_1_onLanes_0_doIt;
  reg                 TrapPlugin_logic_harts_0_crsPorts_write_valid;
  wire                TrapPlugin_logic_harts_0_crsPorts_write_ready;
  reg        [3:0]    TrapPlugin_logic_harts_0_crsPorts_write_address;
  reg        [31:0]   TrapPlugin_logic_harts_0_crsPorts_write_data;
  wire                LsuL1Plugin_logic_bus_read_cmd_valid;
  wire                LsuL1Plugin_logic_bus_read_cmd_ready;
  wire       [31:0]   LsuL1Plugin_logic_bus_read_cmd_payload_address;
  wire                LsuL1Plugin_logic_bus_read_rsp_valid;
  wire                LsuL1Plugin_logic_bus_read_rsp_ready;
  wire       [63:0]   LsuL1Plugin_logic_bus_read_rsp_payload_data;
  wire                LsuL1Plugin_logic_bus_read_rsp_payload_error;
  wire                LsuL1Plugin_logic_bus_write_cmd_valid;
  wire                LsuL1Plugin_logic_bus_write_cmd_ready;
  wire                LsuL1Plugin_logic_bus_write_cmd_payload_last;
  wire       [31:0]   LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address;
  wire       [63:0]   LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data;
  wire                LsuL1Plugin_logic_bus_write_rsp_valid;
  wire                LsuL1Plugin_logic_bus_write_rsp_payload_error;
  reg        [0:0]    LsuL1Plugin_logic_refillCompletions;
  wire                LsuL1Plugin_logic_writebackBusy;
  reg        [3:0]    LsuL1Plugin_logic_banksWrite_mask;
  reg        [8:0]    LsuL1Plugin_logic_banksWrite_address;
  reg        [63:0]   LsuL1Plugin_logic_banksWrite_writeData;
  reg        [7:0]    LsuL1Plugin_logic_banksWrite_writeMask;
  reg        [3:0]    LsuL1Plugin_logic_waysWrite_mask;
  reg        [5:0]    LsuL1Plugin_logic_waysWrite_address;
  reg                 LsuL1Plugin_logic_waysWrite_tag_loaded;
  reg        [19:0]   LsuL1Plugin_logic_waysWrite_tag_address;
  reg                 LsuL1Plugin_logic_waysWrite_tag_fault;
  wire                LsuL1Plugin_logic_waysWrite_valid;
  wire                LsuL1Plugin_logic_banks_0_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_0_write_valid;
  wire       [8:0]    LsuL1Plugin_logic_banks_0_write_payload_address;
  wire       [63:0]   LsuL1Plugin_logic_banks_0_write_payload_data;
  wire       [7:0]    LsuL1Plugin_logic_banks_0_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_0_read_cmd_valid;
  reg        [8:0]    LsuL1Plugin_logic_banks_0_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   LsuL1Plugin_logic_banks_0_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_banks_1_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_1_write_valid;
  wire       [8:0]    LsuL1Plugin_logic_banks_1_write_payload_address;
  wire       [63:0]   LsuL1Plugin_logic_banks_1_write_payload_data;
  wire       [7:0]    LsuL1Plugin_logic_banks_1_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_1_read_cmd_valid;
  reg        [8:0]    LsuL1Plugin_logic_banks_1_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   LsuL1Plugin_logic_banks_1_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_banks_2_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_2_write_valid;
  wire       [8:0]    LsuL1Plugin_logic_banks_2_write_payload_address;
  wire       [63:0]   LsuL1Plugin_logic_banks_2_write_payload_data;
  wire       [7:0]    LsuL1Plugin_logic_banks_2_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_2_read_cmd_valid;
  reg        [8:0]    LsuL1Plugin_logic_banks_2_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   LsuL1Plugin_logic_banks_2_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_banks_3_usedByWriteback;
  wire                LsuL1Plugin_logic_banks_3_write_valid;
  wire       [8:0]    LsuL1Plugin_logic_banks_3_write_payload_address;
  wire       [63:0]   LsuL1Plugin_logic_banks_3_write_payload_data;
  wire       [7:0]    LsuL1Plugin_logic_banks_3_write_payload_mask;
  reg                 LsuL1Plugin_logic_banks_3_read_cmd_valid;
  reg        [8:0]    LsuL1Plugin_logic_banks_3_read_cmd_payload;
  (* keep , syn_keep *) wire       [63:0]   LsuL1Plugin_logic_banks_3_read_rsp /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_0_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded;
  wire                LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_1_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded;
  wire                LsuL1Plugin_logic_ways_2_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_2_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_2_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_2_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_2_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_2_lsuRead_rsp_loaded;
  wire                LsuL1Plugin_logic_ways_3_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_ways_3_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_3_lsuRead_rsp_loaded /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [19:0]   LsuL1Plugin_logic_ways_3_lsuRead_rsp_address /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire                LsuL1Plugin_logic_ways_3_lsuRead_rsp_fault /* synthesis syn_keep = 1 */ ;
  wire       [21:0]   _zz_LsuL1Plugin_logic_ways_3_lsuRead_rsp_loaded;
  reg                 LsuL1Plugin_logic_shared_write_valid;
  reg        [5:0]    LsuL1Plugin_logic_shared_write_payload_address;
  reg        [0:0]    LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  reg        [1:0]    LsuL1Plugin_logic_shared_write_payload_data_plru_1;
  reg        [3:0]    LsuL1Plugin_logic_shared_write_payload_data_dirty;
  wire                LsuL1Plugin_logic_shared_lsuRead_cmd_valid;
  wire       [5:0]    LsuL1Plugin_logic_shared_lsuRead_cmd_payload;
  (* keep , syn_keep *) wire       [0:0]    LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [1:0]    LsuL1Plugin_logic_shared_lsuRead_rsp_plru_1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [3:0]    LsuL1Plugin_logic_shared_lsuRead_rsp_dirty /* synthesis syn_keep = 1 */ ;
  wire       [6:0]    _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_dirty;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0;
  reg                 LsuL1Plugin_logic_refill_slots_0_valid;
  reg                 LsuL1Plugin_logic_refill_slots_0_dirty;
  reg        [31:0]   LsuL1Plugin_logic_refill_slots_0_address;
  reg        [1:0]    LsuL1Plugin_logic_refill_slots_0_way;
  reg                 LsuL1Plugin_logic_refill_slots_0_cmdSent;
  reg                 LsuL1Plugin_logic_refill_slots_0_loadedSet;
  reg                 LsuL1Plugin_logic_refill_slots_0_loaded;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_loadedCounter;
  wire                LsuL1Plugin_logic_refill_slots_0_loadedDone;
  wire                LsuL1Plugin_logic_refill_slots_0_free;
  wire                LsuL1Plugin_logic_refill_slots_0_fire;
  reg        [0:0]    LsuL1Plugin_logic_refill_slots_0_victim;
  wire       [0:0]    LsuL1Plugin_logic_refill_free;
  wire                LsuL1Plugin_logic_refill_full;
  reg                 LsuL1Plugin_logic_refill_push_valid;
  wire       [31:0]   LsuL1Plugin_logic_refill_push_payload_address;
  reg        [1:0]    LsuL1Plugin_logic_refill_push_payload_way;
  reg        [0:0]    LsuL1Plugin_logic_refill_push_payload_victim;
  wire                LsuL1Plugin_logic_refill_push_payload_dirty;
  wire                LsuL1Plugin_logic_refill_push_payload_unique;
  wire                LsuL1Plugin_logic_refill_push_payload_data;
  reg        [31:0]   LsuL1Plugin_logic_refill_pushCounter;
  wire                when_LsuL1Plugin_l377;
  wire                when_LsuL1Plugin_l381;
  wire                LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0;
  wire       [0:0]    LsuL1Plugin_logic_refill_read_arbiter_hits;
  wire                LsuL1Plugin_logic_refill_read_arbiter_hit;
  reg        [0:0]    LsuL1Plugin_logic_refill_read_arbiter_oh;
  reg        [0:0]    LsuL1Plugin_logic_refill_read_arbiter_lock;
  wire                when_LsuL1Plugin_l301;
  wire                LsuL1Plugin_logic_bus_read_cmd_fire;
  wire       [31:0]   LsuL1Plugin_logic_refill_read_cmdAddress;
  wire       [31:0]   LsuL1Plugin_logic_refill_read_rspAddress;
  wire                LsuL1Plugin_logic_refill_read_dirty;
  wire       [1:0]    LsuL1Plugin_logic_refill_read_way;
  (* keep , syn_keep *) reg        [2:0]    LsuL1Plugin_logic_refill_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_refill_read_rspWithData;
  reg        [3:0]    LsuL1Plugin_logic_refill_read_bankWriteNotif;
  wire                LsuL1Plugin_logic_refill_read_writeReservation_win;
  reg                 LsuL1Plugin_logic_refill_read_writeReservation_take;
  reg                 LsuL1Plugin_logic_refill_read_hadError;
  wire                when_LsuL1Plugin_l450;
  reg                 LsuL1Plugin_logic_refill_read_fire;
  wire                LsuL1Plugin_logic_refill_read_reservation_win;
  reg                 LsuL1Plugin_logic_refill_read_reservation_take;
  wire                LsuL1Plugin_logic_refill_read_faulty;
  wire                when_LsuL1Plugin_l463;
  wire       [0:0]    LsuL1_REFILL_BUSY;
  reg                 LsuL1Plugin_logic_writeback_slots_0_fire;
  reg                 LsuL1Plugin_logic_writeback_slots_0_valid;
  reg                 LsuL1Plugin_logic_writeback_slots_0_busy;
  reg        [31:0]   LsuL1Plugin_logic_writeback_slots_0_address;
  reg        [1:0]    LsuL1Plugin_logic_writeback_slots_0_way;
  reg                 LsuL1Plugin_logic_writeback_slots_0_readCmdDone;
  reg                 LsuL1Plugin_logic_writeback_slots_0_readRspDone;
  reg                 LsuL1Plugin_logic_writeback_slots_0_victimBufferReady;
  reg                 LsuL1Plugin_logic_writeback_slots_0_writeCmdDone;
  reg        [0:0]    LsuL1Plugin_logic_writeback_slots_0_timer_counter;
  wire                LsuL1Plugin_logic_writeback_slots_0_timer_done;
  wire                when_LsuL1Plugin_l530;
  wire                LsuL1Plugin_logic_writeback_slots_0_free;
  wire       [0:0]    LsuL1_WRITEBACK_BUSY;
  wire       [0:0]    LsuL1Plugin_logic_writeback_free;
  wire                LsuL1Plugin_logic_writeback_full;
  reg                 LsuL1Plugin_logic_writeback_push_valid;
  reg        [31:0]   LsuL1Plugin_logic_writeback_push_payload_address;
  reg        [1:0]    LsuL1Plugin_logic_writeback_push_payload_way;
  wire                when_LsuL1Plugin_l556;
  wire                when_LsuL1Plugin_l561;
  wire                LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0;
  wire       [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_hits;
  wire                LsuL1Plugin_logic_writeback_read_arbiter_hit;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_oh;
  reg        [0:0]    LsuL1Plugin_logic_writeback_read_arbiter_lock;
  wire                when_LsuL1Plugin_l301_1;
  wire       [31:0]   LsuL1Plugin_logic_writeback_read_address;
  wire       [1:0]    LsuL1Plugin_logic_writeback_read_way;
  (* keep , syn_keep *) reg        [2:0]    LsuL1Plugin_logic_writeback_read_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_writeback_read_slotRead_valid;
  wire                LsuL1Plugin_logic_writeback_read_slotRead_payload_last;
  wire       [2:0]    LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex;
  wire       [1:0]    LsuL1Plugin_logic_writeback_read_slotRead_payload_way;
  wire                when_LsuL1Plugin_l605;
  reg                 LsuL1Plugin_logic_writeback_read_slotReadLast_valid;
  reg                 LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last;
  reg        [2:0]    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex;
  reg        [1:0]    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way;
  wire       [63:0]   LsuL1Plugin_logic_writeback_read_readedData;
  wire                LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0;
  wire       [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_hits;
  wire                LsuL1Plugin_logic_writeback_write_arbiter_hit;
  reg        [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_oh;
  reg        [0:0]    LsuL1Plugin_logic_writeback_write_arbiter_lock;
  wire                when_LsuL1Plugin_l301_2;
  (* keep , syn_keep *) reg        [2:0]    LsuL1Plugin_logic_writeback_write_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                LsuL1Plugin_logic_writeback_write_last;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_valid;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_ready;
  wire       [31:0]   LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_payload_last;
  wire                LsuL1Plugin_logic_writeback_write_bufferRead_fire;
  wire                when_LsuL1Plugin_l676;
  wire                LsuL1Plugin_logic_writeback_write_cmd_valid;
  wire                LsuL1Plugin_logic_writeback_write_cmd_ready;
  wire       [31:0]   LsuL1Plugin_logic_writeback_write_cmd_payload_address;
  wire                LsuL1Plugin_logic_writeback_write_cmd_payload_last;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_rValid;
  reg        [31:0]   LsuL1Plugin_logic_writeback_write_bufferRead_rData_address;
  reg                 LsuL1Plugin_logic_writeback_write_bufferRead_rData_last;
  wire                when_Stream_l399;
  wire       [2:0]    _zz_LsuL1Plugin_logic_writeback_write_word;
  wire       [63:0]   LsuL1Plugin_logic_writeback_write_word;
  wire       [8:0]    LsuL1Plugin_logic_lsu_rb0_readAddress;
  wire                when_LsuL1Plugin_l718;
  wire                when_LsuL1Plugin_l719;
  wire                when_LsuL1Plugin_l718_1;
  wire                when_LsuL1Plugin_l719_1;
  wire                when_LsuL1Plugin_l718_2;
  wire                when_LsuL1Plugin_l719_2;
  wire                when_LsuL1Plugin_l718_3;
  wire                when_LsuL1Plugin_l719_3;
  reg                 LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg;
  wire                when_LsuL1Plugin_l735;
  reg                 LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg;
  wire                when_LsuL1Plugin_l735_1;
  reg                 LsuL1Plugin_logic_lsu_rb1_onBanks_2_busyReg;
  wire                when_LsuL1Plugin_l735_2;
  reg                 LsuL1Plugin_logic_lsu_rb1_onBanks_3_busyReg;
  wire                when_LsuL1Plugin_l735_3;
  wire                _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
  wire                _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1;
  wire                _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_2;
  wire                _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_3;
  wire                LsuL1Plugin_logic_lsu_sharedBypassers_0_hit;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_0;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_1;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_evict_id;
  reg        [1:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_0;
  reg        [1:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_1;
  wire                LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_1;
  wire                LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_0_state;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_1_stateSel;
  wire                LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_1_state;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_update_logic_1_sel;
  wire                LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win;
  reg                 LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take;
  wire                LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win;
  wire                LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_take;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate;
  wire                LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_refillHazards;
  wire       [0:0]    LsuL1Plugin_logic_lsu_ctrl_writebackHazards;
  wire                LsuL1Plugin_logic_lsu_ctrl_refillHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_writebackHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_wasDirty;
  wire       [3:0]    LsuL1Plugin_logic_lsu_ctrl_loadedDirties;
  wire                LsuL1Plugin_logic_lsu_ctrl_refillWayWasDirty;
  wire                LsuL1Plugin_logic_lsu_ctrl_writeToReadHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_bankNotRead;
  wire                LsuL1Plugin_logic_lsu_ctrl_loadHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_storeHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_preventSideEffects;
  wire                LsuL1Plugin_logic_lsu_ctrl_flushHazard;
  wire                LsuL1Plugin_logic_lsu_ctrl_coherencyHazard;
  reg                 LsuL1Plugin_logic_lsu_ctrl_hazardReg;
  reg                 LsuL1Plugin_logic_lsu_ctrl_flushHazardReg;
  wire                LsuL1Plugin_logic_lsu_ctrl_canRefill;
  wire                LsuL1Plugin_logic_lsu_ctrl_canFlush;
  wire       [3:0]    LsuL1Plugin_logic_lsu_ctrl_needFlushs;
  wire       [3:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_2;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_3;
  reg        [3:0]    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_range_0_to_1;
  wire                LsuL1Plugin_logic_lsu_ctrl_needFlushs_range_0_to_2;
  wire       [3:0]    LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
  wire                _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
  wire                _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel_1;
  wire                _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel_2;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
  wire                LsuL1Plugin_logic_lsu_ctrl_isAccess;
  wire                LsuL1Plugin_logic_lsu_ctrl_askRefill;
  wire                LsuL1Plugin_logic_lsu_ctrl_askUpgrade;
  wire                LsuL1Plugin_logic_lsu_ctrl_askFlush;
  wire                LsuL1Plugin_logic_lsu_ctrl_askCbm;
  wire                LsuL1Plugin_logic_lsu_ctrl_doRefill;
  wire                LsuL1Plugin_logic_lsu_ctrl_doUpgrade;
  wire                LsuL1Plugin_logic_lsu_ctrl_doFlush;
  wire                LsuL1Plugin_logic_lsu_ctrl_doWrite;
  wire                LsuL1Plugin_logic_lsu_ctrl_doCbm;
  wire                _zz_LsuL1Plugin_logic_lsu_ctrl_wayId;
  wire                _zz_LsuL1Plugin_logic_lsu_ctrl_wayId_1;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_wayId;
  wire       [1:0]    LsuL1Plugin_logic_lsu_ctrl_targetWay;
  wire       [2:0]    _zz_45;
  wire       [2:0]    _zz_46;
  wire       [2:0]    _zz_47;
  wire       [2:0]    _zz_48;
  wire       [2:0]    _zz_49;
  wire       [2:0]    _zz_50;
  wire       [2:0]    _zz_51;
  wire       [2:0]    _zz_52;
  wire                LsuL1Plugin_logic_lsu_ctrl_doRefillPush;
  wire                when_LsuL1Plugin_l915;
  wire       [2:0]    _zz_53;
  wire       [1:0]    _zz_54;
  wire                when_LsuL1Plugin_l929;
  wire                when_LsuL1Plugin_l929_1;
  wire                when_LsuL1Plugin_l929_2;
  wire                when_LsuL1Plugin_l929_3;
  wire       [19:0]   _zz_LsuL1Plugin_logic_waysWrite_tag_address;
  wire                when_LsuL1Plugin_l1019;
  wire                when_LsuL1Plugin_l1026;
  wire                when_LsuL1Plugin_l1030;
  wire                when_LsuL1Plugin_l1030_1;
  wire                when_LsuL1Plugin_l1030_2;
  wire                when_LsuL1Plugin_l1030_3;
  wire                when_LsuL1Plugin_l1026_1;
  wire                when_LsuL1Plugin_l1030_4;
  wire                when_LsuL1Plugin_l1030_5;
  wire                when_LsuL1Plugin_l1030_6;
  wire                when_LsuL1Plugin_l1030_7;
  reg        [6:0]    LsuL1Plugin_logic_initializer_counter;
  wire                LsuL1Plugin_logic_initializer_done;
  wire                when_LsuL1Plugin_l1219;
  wire       [6:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty;
  wire       [2:0]    _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  reg                 TrapPlugin_logic_harts_0_interrupt_valid;
  reg        [3:0]    TrapPlugin_logic_harts_0_interrupt_code;
  reg        [1:0]    TrapPlugin_logic_harts_0_interrupt_targetPrivilege;
  wire                when_TrapPlugin_l201;
  wire                when_TrapPlugin_l201_1;
  wire                when_TrapPlugin_l207;
  wire                when_TrapPlugin_l207_1;
  wire                when_TrapPlugin_l207_2;
  wire                when_TrapPlugin_l207_3;
  wire                when_TrapPlugin_l207_4;
  wire                when_TrapPlugin_l207_5;
  wire                when_TrapPlugin_l207_6;
  wire                when_TrapPlugin_l207_7;
  wire                when_TrapPlugin_l207_8;
  reg                 TrapPlugin_logic_harts_0_interrupt_validBuffer;
  wire                TrapPlugin_logic_harts_0_interrupt_pendingInterrupt;
  wire                when_TrapPlugin_l226;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg;
  wire       [1:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception;
  wire       [39:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_arg;
  wire       [4:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3;
  wire                _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4;
  reg        [4:0]    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_5;
  wire       [4:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_oh;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid;
  wire                TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code;
  wire       [2:0]    TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg;
  wire       [39:0]   _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
  reg                 TrapPlugin_logic_harts_0_trap_pending_state_exception;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_pending_state_tval;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_pending_state_code;
  reg        [2:0]    TrapPlugin_logic_harts_0_trap_pending_state_arg;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_pending_pc;
  reg        [11:0]   TrapPlugin_logic_harts_0_trap_pending_history;
  reg        [0:0]    TrapPlugin_logic_harts_0_trap_pending_slices;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_exception_code;
  wire                when_TrapPlugin_l263;
  wire                when_TrapPlugin_l263_1;
  wire                when_TrapPlugin_l263_2;
  wire                when_TrapPlugin_l263_3;
  wire                when_TrapPlugin_l263_4;
  wire                when_TrapPlugin_l263_5;
  wire                when_TrapPlugin_l263_6;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_exception_targetPrivilege;
  wire                execute_lane0_ctrls_5_upIsCancel;
  wire                execute_lane0_ctrls_5_downIsCancel;
  wire       [0:0]    TrapPlugin_logic_harts_0_trap_trigger_oh;
  wire                TrapPlugin_logic_harts_0_trap_trigger_valid;
  reg                 TrapPlugin_logic_harts_0_trap_whitebox_trap;
  reg                 TrapPlugin_logic_harts_0_trap_whitebox_interrupt;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_whitebox_code;
  reg                 TrapPlugin_logic_harts_0_trap_historyPort_valid;
  wire       [11:0]   TrapPlugin_logic_harts_0_trap_historyPort_payload_history;
  reg                 TrapPlugin_logic_harts_0_trap_pcPort_valid;
  wire                TrapPlugin_logic_harts_0_trap_pcPort_payload_fault;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_pcPort_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_wantExit;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_wantStart;
  wire                TrapPlugin_logic_harts_0_trap_fsm_wantKill;
  wire                TrapPlugin_logic_harts_0_trap_fsm_inflightTrap;
  wire                TrapPlugin_logic_harts_0_trap_fsm_holdPort;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_wfi;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code;
  reg        [1:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege;
  wire                TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval;
  wire       [3:0]    TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
  wire                TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_ready;
  wire       [31:0]   TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_address;
  wire       [0:0]    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_storageId;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid;
  wire                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated;
  wire                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_fire;
  wire                when_TrapPlugin_l355;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
  wire       [0:0]    TrapPlugin_logic_harts_0_trap_fsm_jumpOffset;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug;
  wire                TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak;
  reg                 TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg;
  wire                when_TrapPlugin_l556;
  reg        [31:0]   TrapPlugin_logic_harts_0_trap_fsm_readed;
  wire       [1:0]    TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege;
  reg        [0:0]    LsuPlugin_logic_flusher_waiter;
  wire       [4:0]    LsuPlugin_logic_onAddress0_ls_prefetchOp;
  wire                LsuPlugin_logic_onAddress0_ls_port_valid;
  wire                LsuPlugin_logic_onAddress0_ls_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_ls_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_ls_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_ls_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_ls_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_ls_port_payload_storeId;
  reg        [11:0]   LsuPlugin_logic_onAddress0_ls_storeId;
  wire                LsuPlugin_logic_onAddress0_ls_port_fire;
  reg        [0:0]    LsuPlugin_logic_onAddress0_access_waiter_refill;
  reg                 LsuPlugin_logic_onAddress0_access_waiter_valid;
  wire                when_LsuPlugin_l259;
  wire                LsuPlugin_logic_onAddress0_access_sbWaiter;
  wire                LsuPlugin_logic_onAddress0_access_port_valid;
  wire                LsuPlugin_logic_onAddress0_access_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_access_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_access_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_access_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_access_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_access_port_payload_storeId;
  wire                _zz_MmuPlugin_logic_accessBus_cmd_ready;
  wire                MmuPlugin_logic_accessBus_cmd_haltWhen_valid;
  wire                MmuPlugin_logic_accessBus_cmd_haltWhen_ready;
  wire       [31:0]   MmuPlugin_logic_accessBus_cmd_haltWhen_payload_address;
  wire       [1:0]    MmuPlugin_logic_accessBus_cmd_haltWhen_payload_size;
  wire                LsuPlugin_logic_onAddress0_flush_port_valid;
  wire                LsuPlugin_logic_onAddress0_flush_port_ready;
  wire       [2:0]    LsuPlugin_logic_onAddress0_flush_port_payload_op;
  wire       [31:0]   LsuPlugin_logic_onAddress0_flush_port_payload_address;
  wire       [1:0]    LsuPlugin_logic_onAddress0_flush_port_payload_size;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_load;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_store;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_atomic;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_clean;
  wire                LsuPlugin_logic_onAddress0_flush_port_payload_invalidate;
  wire       [11:0]   LsuPlugin_logic_onAddress0_flush_port_payload_storeId;
  wire                LsuPlugin_logic_onAddress0_flush_port_fire;
  reg        [3:0]    _zz_execute_ctrl2_down_LsuL1_MASK_lane0;
  wire                when_LsuPlugin_l546;
  wire                when_LsuPlugin_l546_1;
  wire       [31:0]   LsuPlugin_logic_onPma_cached_cmd_address;
  wire       [0:0]    LsuPlugin_logic_onPma_cached_cmd_op;
  wire                LsuPlugin_logic_onPma_cached_rsp_fault;
  wire                LsuPlugin_logic_onPma_cached_rsp_io;
  wire       [31:0]   LsuPlugin_logic_onPma_io_cmd_address;
  wire       [1:0]    LsuPlugin_logic_onPma_io_cmd_size;
  wire       [0:0]    LsuPlugin_logic_onPma_io_cmd_op;
  wire                LsuPlugin_logic_onPma_io_rsp_fault;
  wire                LsuPlugin_logic_onPma_io_rsp_io;
  wire                when_LsuPlugin_l569;
  wire                LsuPlugin_logic_onPma_addressExtension;
  reg                 LsuPlugin_logic_onCtrl_lsuTrap;
  reg        [31:0]   LsuPlugin_logic_onCtrl_writeData;
  wire                LsuPlugin_logic_onCtrl_scMiss;
  reg                 LsuPlugin_logic_onCtrl_io_tooEarly;
  reg                 LsuPlugin_logic_onCtrl_io_allowIt;
  wire                when_LsuPlugin_l597;
  wire                LsuPlugin_logic_onCtrl_io_doIt;
  reg                 LsuPlugin_logic_onCtrl_io_doItReg;
  reg                 LsuPlugin_logic_onCtrl_io_cmdSent;
  wire                LsuPlugin_logic_bus_cmd_fire;
  wire                when_LsuPlugin_l601;
  wire                LsuPlugin_logic_bus_rsp_toStream_valid;
  wire                LsuPlugin_logic_bus_rsp_toStream_ready;
  wire                LsuPlugin_logic_bus_rsp_toStream_payload_error;
  wire       [31:0]   LsuPlugin_logic_bus_rsp_toStream_payload_data;
  wire                LsuPlugin_logic_onCtrl_io_rsp_valid;
  wire                LsuPlugin_logic_onCtrl_io_rsp_ready;
  wire                LsuPlugin_logic_onCtrl_io_rsp_payload_error;
  wire       [31:0]   LsuPlugin_logic_onCtrl_io_rsp_payload_data;
  reg                 LsuPlugin_logic_bus_rsp_toStream_rValid;
  wire                LsuPlugin_logic_onCtrl_io_rsp_fire;
  reg                 LsuPlugin_logic_bus_rsp_toStream_rData_error;
  reg        [31:0]   LsuPlugin_logic_bus_rsp_toStream_rData_data;
  wire                LsuPlugin_logic_onCtrl_io_freezeIt;
  wire       [31:0]   LsuPlugin_logic_onCtrl_loadData_input;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_0;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_1;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_2;
  wire       [7:0]    LsuPlugin_logic_onCtrl_loadData_splitted_3;
  reg        [31:0]   LsuPlugin_logic_onCtrl_loadData_shifted;
  wire       [31:0]   LsuPlugin_logic_onCtrl_storeData_mapping_0_1;
  wire       [31:0]   LsuPlugin_logic_onCtrl_storeData_mapping_1_1;
  wire       [31:0]   LsuPlugin_logic_onCtrl_storeData_mapping_2_1;
  reg        [31:0]   _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_srcBuffer;
  wire       [2:0]    _zz_LsuPlugin_logic_onCtrl_rva_alu_compare;
  wire                _zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf;
  wire                LsuPlugin_logic_onCtrl_rva_alu_compare;
  wire                LsuPlugin_logic_onCtrl_rva_alu_unsigned;
  wire       [31:0]   LsuPlugin_logic_onCtrl_rva_alu_addSub;
  wire                LsuPlugin_logic_onCtrl_rva_alu_less;
  wire                LsuPlugin_logic_onCtrl_rva_alu_selectRf;
  wire       [2:0]    switch_Misc_l242_1;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_alu_raw;
  wire       [31:0]   LsuPlugin_logic_onCtrl_rva_alu_result;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_aluBuffer;
  wire                LsuPlugin_logic_onCtrl_rva_delay_0;
  wire                LsuPlugin_logic_onCtrl_rva_delay_1;
  reg                 _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
  reg                 _zz_LsuPlugin_logic_onCtrl_rva_delay_1;
  wire                LsuPlugin_logic_onCtrl_rva_freezeIt;
  reg                 LsuPlugin_logic_onCtrl_rva_lrsc_capture;
  reg                 LsuPlugin_logic_onCtrl_rva_lrsc_reserved;
  reg        [31:0]   LsuPlugin_logic_onCtrl_rva_lrsc_address;
  wire                when_LsuPlugin_l685;
  reg        [5:0]    LsuPlugin_logic_onCtrl_rva_lrsc_age;
  wire                when_LsuPlugin_l697;
  wire                LsuPlugin_logic_onCtrl_traps_accessFault;
  wire                LsuPlugin_logic_onCtrl_traps_l1Failed;
  wire                LsuPlugin_logic_onCtrl_traps_pmaFault;
  wire                when_LsuPlugin_l806;
  wire                when_LsuPlugin_l833;
  wire                when_LsuPlugin_l861;
  wire                LsuPlugin_logic_onCtrl_mmuNeeded;
  wire                when_LsuPlugin_l901;
  wire                when_LsuPlugin_l938;
  wire                when_LsuPlugin_l263;
  reg        [0:0]    LsuPlugin_logic_onCtrl_hartRegulation_refill;
  reg                 LsuPlugin_logic_onCtrl_hartRegulation_valid;
  wire                when_LsuPlugin_l259_1;
  wire                when_LsuPlugin_l945;
  wire                when_LsuPlugin_l263_1;
  wire                when_LsuPlugin_l968;
  wire                LsuPlugin_logic_onWb_storeFire;
  wire                LsuPlugin_logic_onWb_storeBroadcast;
  reg                 LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock;
  wire                LsuL1TileLinkPlugin_logic_down_a_fire;
  reg        [2:0]    LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat;
  wire                LsuL1TileLinkPlugin_logic_down_a_tracker_last;
  wire                when_LsuL1Bus_l151;
  reg                 LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_selReg;
  wire                LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel;
  wire                LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel;
  wire                PcPlugin_logic_forcedSpawn;
  reg        [9:0]    PcPlugin_logic_harts_0_self_id;
  wire                PcPlugin_logic_harts_0_self_flow_valid;
  wire                PcPlugin_logic_harts_0_self_flow_payload_fault;
  wire       [31:0]   PcPlugin_logic_harts_0_self_flow_payload_pc;
  wire                PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid;
  reg                 PcPlugin_logic_harts_0_self_increment;
  reg                 PcPlugin_logic_harts_0_self_fault;
  reg        [31:0]   PcPlugin_logic_harts_0_self_state;
  wire       [31:0]   PcPlugin_logic_harts_0_self_pc;
  wire                PcPlugin_logic_harts_0_aggregator_valids_0;
  wire                PcPlugin_logic_harts_0_aggregator_valids_1;
  wire                PcPlugin_logic_harts_0_aggregator_valids_2;
  wire                PcPlugin_logic_harts_0_aggregator_valids_3;
  wire       [3:0]    _zz_PcPlugin_logic_harts_0_aggregator_oh;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_1;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_2;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_oh_3;
  reg        [3:0]    _zz_PcPlugin_logic_harts_0_aggregator_oh_4;
  wire       [3:0]    PcPlugin_logic_harts_0_aggregator_oh;
  (* keep , syn_keep *) wire       [31:0]   PcPlugin_logic_harts_0_aggregator_target /* synthesis syn_keep = 1 */ ;
  wire                PcPlugin_logic_harts_0_aggregator_fault;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_1;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_target_2;
  wire                _zz_PcPlugin_logic_harts_0_aggregator_fault_1;
  wire                when_PcPlugin_l80;
  wire                PcPlugin_logic_harts_0_holdComb;
  reg                 PcPlugin_logic_harts_0_holdReg;
  wire                PcPlugin_logic_harts_0_output_valid;
  wire                PcPlugin_logic_harts_0_output_ready;
  reg        [31:0]   PcPlugin_logic_harts_0_output_payload_pc;
  wire                PcPlugin_logic_harts_0_output_payload_fault;
  wire                PcPlugin_logic_harts_0_output_fire;
  wire                PcPlugin_logic_holdHalter_doIt;
  wire                fetch_logic_ctrls_0_haltRequest_PcPlugin_l133;
  reg        [11:0]   HistoryPlugin_logic_onFetch_value;
  reg        [11:0]   HistoryPlugin_logic_onFetch_valueNext;
  wire                HistoryPlugin_logic_onFetch_ports_0_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_0_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_1_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_1_payload_history;
  wire                HistoryPlugin_logic_onFetch_ports_2_valid;
  wire       [11:0]   HistoryPlugin_logic_onFetch_ports_2_payload_history;
  reg        [1:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask;
  reg        [4:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid;
  reg        [14:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willClear;
  reg        [0:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [0:0]    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [0:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask;
  reg        [4:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid;
  reg        [4:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [9:0]    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willClear;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflow;
  reg        [2:0]    LsuPlugin_logic_translationStorage_logic_sl_0_write_mask;
  reg        [4:0]    LsuPlugin_logic_translationStorage_logic_sl_0_write_address;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid;
  reg        [14:0]   LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress;
  reg        [19:0]   LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willClear;
  reg        [1:0]    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
  reg        [1:0]    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc;
  wire                LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflow;
  reg        [0:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_mask;
  reg        [4:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_address;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid;
  reg        [4:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress;
  reg        [9:0]    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser;
  reg                 LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willClear;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc;
  wire                LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflow;
  wire                MmuPlugin_logic_isMachine;
  wire                MmuPlugin_logic_isSupervisor;
  wire                MmuPlugin_logic_isUser;
  wire                when_MmuPlugin_l275;
  wire                when_MmuPlugin_l277;
  wire       [4:0]    LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress;
  wire       [39:0]   _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid;
  wire       [39:0]   _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid;
  wire       [39:0]   _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid;
  wire       [4:0]    LsuPlugin_logic_onAddress0_translationPort_logic_read_1_readAddress;
  wire       [19:0]   _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid;
  wire       [3:0]    LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hit;
  wire       [3:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_3;
  reg        [3:0]    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_1;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_2;
  wire       [3:0]    LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite;
  wire                LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser;
  wire       [31:0]   LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated;
  reg                 LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup;
  wire       [4:0]    FetchL1Plugin_logic_translationPort_logic_read_0_readAddress;
  wire       [39:0]   _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid;
  wire       [39:0]   _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid;
  wire       [4:0]    FetchL1Plugin_logic_translationPort_logic_read_1_readAddress;
  wire       [19:0]   _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid;
  wire       [2:0]    FetchL1Plugin_logic_translationPort_logic_ctrl_hits;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hit;
  wire       [2:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_2;
  reg        [2:0]    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_hits_range_0_to_1;
  wire       [2:0]    FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  wire                _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1;
  wire                _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite;
  wire                FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser;
  wire       [31:0]   FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated;
  reg                 FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup;
  wire                MmuPlugin_logic_refill_wantExit;
  reg                 MmuPlugin_logic_refill_wantStart;
  wire                MmuPlugin_logic_refill_wantKill;
  wire                MmuPlugin_logic_refill_busy;
  reg        [31:0]   MmuPlugin_logic_refill_virtual;
  reg                 MmuPlugin_logic_refill_cacheRefillAny;
  reg                 MmuPlugin_logic_refill_cacheRefillAnySet;
  reg        [0:0]    MmuPlugin_logic_refill_portOhReg;
  reg        [1:0]    MmuPlugin_logic_refill_storageOhReg;
  wire                MmuPlugin_logic_refill_events_onStorage_0_waiting;
  wire                MmuPlugin_logic_refill_events_onStorage_1_waiting;
  reg        [31:0]   MmuPlugin_logic_refill_load_address;
  reg                 MmuPlugin_logic_refill_load_rsp_valid;
  reg        [31:0]   MmuPlugin_logic_refill_load_rsp_payload_data;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_error;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_redo;
  reg                 MmuPlugin_logic_refill_load_rsp_payload_waitAny;
  wire       [31:0]   MmuPlugin_logic_refill_load_readed;
  wire                when_MmuPlugin_l395;
  wire                MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_flags_R;
  wire                MmuPlugin_logic_refill_load_flags_W;
  wire                MmuPlugin_logic_refill_load_flags_X;
  wire                MmuPlugin_logic_refill_load_flags_U;
  wire                MmuPlugin_logic_refill_load_flags_G;
  wire                MmuPlugin_logic_refill_load_flags_A;
  wire                MmuPlugin_logic_refill_load_flags_D;
  wire       [31:0]   _zz_MmuPlugin_logic_refill_load_flags_V;
  wire                MmuPlugin_logic_refill_load_leaf;
  wire                MmuPlugin_logic_refill_load_reservedFault;
  reg                 MmuPlugin_logic_refill_load_exception;
  reg        [31:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_0;
  reg        [31:0]   MmuPlugin_logic_refill_load_levelToPhysicalAddress_1;
  wire                MmuPlugin_logic_refill_load_levelException_0;
  reg                 MmuPlugin_logic_refill_load_levelException_1;
  reg        [31:0]   MmuPlugin_logic_refill_load_nextLevelBase;
  wire                when_MmuPlugin_l416;
  wire                MmuPlugin_logic_refill_fetch_0_pteFault;
  wire                MmuPlugin_logic_refill_fetch_0_leafAccessFault;
  wire                MmuPlugin_logic_refill_fetch_0_pageFault;
  wire                MmuPlugin_logic_refill_fetch_0_accessFault;
  wire                MmuPlugin_logic_refill_fetch_1_pteFault;
  wire                MmuPlugin_logic_refill_fetch_1_leafAccessFault;
  wire                MmuPlugin_logic_refill_fetch_1_pageFault;
  wire                MmuPlugin_logic_refill_fetch_1_accessFault;
  reg        [4:0]    MmuPlugin_logic_invalidate_counter;
  reg                 MmuPlugin_logic_invalidate_busy;
  wire                when_MmuPlugin_l512;
  wire                when_MmuPlugin_l526;
  wire                PmpPlugin_logic_isMachine;
  wire                PmpPlugin_logic_instructionShouldHit;
  wire                PmpPlugin_logic_dataShouldHit;
  wire                FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort;
  wire       [19:0]   FetchL1Plugin_logic_pmpPort_logic_torCmpAddress;
  wire                LsuPlugin_logic_pmpPort_logic_dataShouldHitPort;
  wire       [19:0]   LsuPlugin_logic_pmpPort_logic_torCmpAddress;
  wire       [7:0]    LsuTileLinkPlugin_logic_bridge_cmdHash;
  wire       [2:0]    _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode;
  wire                fetch_logic_flushes_0_doIt;
  wire                fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48;
  wire                fetch_logic_flushes_1_doIt;
  wire                fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l50;
  reg                 PerformanceCounterPlugin_logic_interrupt_ip;
  reg                 PerformanceCounterPlugin_logic_interrupt_ie;
  reg                 PerformanceCounterPlugin_logic_interrupt_sup_deleg;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_0;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_0;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_1;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_1;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_2;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_2;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_3;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_3;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_4;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_4;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_5;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_5;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_6;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_6;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_7;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_7;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_8;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_8;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_9;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_9;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_10;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_10;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_11;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_11;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_12;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_12;
  reg        [0:0]    _zz_PerformanceCounterPlugin_logic_events_sums_13;
  wire       [0:0]    PerformanceCounterPlugin_logic_events_sums_13;
  wire                PerformanceCounterPlugin_logic_fsm_wantExit;
  reg                 PerformanceCounterPlugin_logic_fsm_wantStart;
  wire                PerformanceCounterPlugin_logic_fsm_wantKill;
  wire                PerformanceCounterPlugin_logic_fsm_flusherCmd_valid;
  reg                 PerformanceCounterPlugin_logic_fsm_flusherCmd_ready;
  wire       [1:0]    PerformanceCounterPlugin_logic_fsm_flusherCmd_payload_oh;
  reg                 PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid;
  reg                 PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready;
  wire       [1:0]    PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address;
  wire                PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid;
  reg                 PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready;
  wire       [1:0]    PerformanceCounterPlugin_logic_fsm_csrReadCmd_payload_address;
  reg                 PerformanceCounterPlugin_logic_fsm_cmd_flusher;
  reg        [1:0]    PerformanceCounterPlugin_logic_fsm_cmd_oh;
  wire                _zz_PerformanceCounterPlugin_logic_fsm_cmd_address;
  wire                _zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1;
  wire       [2:0]    PerformanceCounterPlugin_logic_fsm_cmd_address;
  wire                PerformanceCounterPlugin_logic_fsm_done;
  reg        [31:0]   PerformanceCounterPlugin_logic_fsm_ramReaded;
  reg                 PerformanceCounterPlugin_logic_fsm_carry;
  reg        [7:0]    PerformanceCounterPlugin_logic_fsm_counterReaded;
  wire       [31:0]   PerformanceCounterPlugin_logic_fsm_calc_a;
  wire       [7:0]    PerformanceCounterPlugin_logic_fsm_calc_b;
  wire       [32:0]   PerformanceCounterPlugin_logic_fsm_calc_sum;
  wire       [1:0]    PerformanceCounterPlugin_logic_fsm_idleCsrAddress;
  reg                 PerformanceCounterPlugin_logic_fsm_holdCsrWrite;
  wire       [1:0]    PerformanceCounterPlugin_logic_flusher_hits;
  wire                PerformanceCounterPlugin_logic_flusher_hit;
  wire       [1:0]    PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input;
  wire       [1:0]    PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked;
  wire       [1:0]    PerformanceCounterPlugin_logic_flusher_oh;
  wire       [1:0]    PerformanceCounterPlugin_logic_csrDecode_addr;
  reg                 PerformanceCounterPlugin_logic_csrDecode_mok;
  reg                 PerformanceCounterPlugin_logic_csrDecode_sok;
  wire                PerformanceCounterPlugin_logic_csrDecode_privOk;
  reg                 PerformanceCounterPlugin_logic_csrRead_fired;
  wire                PerformanceCounterPlugin_logic_fsm_csrReadCmd_fire;
  wire                PerformanceCounterPlugin_logic_csrRead_requested;
  wire                when_PerformanceCounterPlugin_l342;
  reg                 PerformanceCounterPlugin_logic_csrWrite_fired;
  wire                PerformanceCounterPlugin_logic_fsm_csrWriteCmd_fire;
  wire                CsrAccessPlugin_logic_fsm_wantExit;
  reg                 CsrAccessPlugin_logic_fsm_wantStart;
  wire                CsrAccessPlugin_logic_fsm_wantKill;
  reg                 REG_CSR_768;
  reg                 REG_CSR_256;
  reg                 REG_CSR_384;
  reg                 REG_CSR_3008;
  reg                 REG_CSR_1952;
  reg                 REG_CSR_1953;
  reg                 REG_CSR_1954;
  reg                 REG_CSR_3857;
  reg                 REG_CSR_3858;
  reg                 REG_CSR_3859;
  reg                 REG_CSR_3860;
  reg                 REG_CSR_769;
  reg                 REG_CSR_834;
  reg                 REG_CSR_836;
  reg                 REG_CSR_772;
  reg                 REG_CSR_770;
  reg                 REG_CSR_771;
  reg                 REG_CSR_322;
  reg                 REG_CSR_260;
  reg                 REG_CSR_324;
  reg                 REG_CSR_3073;
  reg                 REG_CSR_3201;
  reg                 REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
  reg                 REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
  reg                 REG_CSR_774;
  reg                 REG_CSR_262;
  reg                 REG_CSR_800;
  reg                 REG_CSR_;
  reg                 REG_CSR_CsrRamPlugin_csrMapper_selFilter;
  reg                 REG_CSR_PerformanceCounterPlugin_logic_csrFilter;
  reg                 REG_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
  reg                 CsrAccessPlugin_logic_fsm_interface_read;
  reg                 CsrAccessPlugin_logic_fsm_interface_write;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_interface_rs1;
  reg        [31:0]   CsrAccessPlugin_logic_fsm_interface_aluInput;
  reg        [31:0]   CsrAccessPlugin_logic_fsm_interface_csrValue;
  reg        [31:0]   CsrAccessPlugin_logic_fsm_interface_onWriteBits;
  wire       [15:0]   CsrAccessPlugin_logic_fsm_interface_uopId;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_interface_uop;
  wire                CsrAccessPlugin_logic_fsm_interface_doImm;
  wire                CsrAccessPlugin_logic_fsm_interface_doMask;
  wire                CsrAccessPlugin_logic_fsm_interface_doClear;
  wire       [4:0]    CsrAccessPlugin_logic_fsm_interface_rdPhys;
  wire                CsrAccessPlugin_logic_fsm_interface_rdEnable;
  reg                 CsrAccessPlugin_logic_fsm_interface_fire;
  wire       [11:0]   CsrAccessPlugin_logic_fsm_inject_csrAddress;
  wire                CsrAccessPlugin_logic_fsm_inject_immZero;
  wire                CsrAccessPlugin_logic_fsm_inject_srcZero;
  wire                CsrAccessPlugin_logic_fsm_inject_csrWrite;
  wire                CsrAccessPlugin_logic_fsm_inject_csrRead;
  wire                COMB_CSR_768;
  wire                COMB_CSR_256;
  wire                COMB_CSR_384;
  wire                COMB_CSR_3008;
  wire                COMB_CSR_1952;
  wire                COMB_CSR_1953;
  wire                COMB_CSR_1954;
  wire                COMB_CSR_3857;
  wire                COMB_CSR_3858;
  wire                COMB_CSR_3859;
  wire                COMB_CSR_3860;
  wire                COMB_CSR_769;
  wire                COMB_CSR_834;
  wire                COMB_CSR_836;
  wire                COMB_CSR_772;
  wire                COMB_CSR_770;
  wire                COMB_CSR_771;
  wire                COMB_CSR_322;
  wire                COMB_CSR_260;
  wire                COMB_CSR_324;
  wire                COMB_CSR_3073;
  wire                COMB_CSR_3201;
  wire                COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
  wire                COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
  wire                COMB_CSR_774;
  wire                COMB_CSR_262;
  wire                COMB_CSR_800;
  wire                COMB_CSR_;
  wire                COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
  wire                COMB_CSR_PerformanceCounterPlugin_logic_csrFilter;
  wire                COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
  wire                CsrAccessPlugin_logic_fsm_inject_implemented;
  wire                CsrAccessPlugin_logic_fsm_inject_onDecodeDo;
  wire                when_CsrAccessPlugin_l155;
  wire                when_MmuPlugin_l221;
  wire                when_CsrAccessPlugin_l155_1;
  wire                when_CsrAccessPlugin_l155_2;
  wire                when_PerformanceCounterPlugin_l327;
  wire                when_PerformanceCounterPlugin_l328;
  wire                when_CsrAccessPlugin_l155_3;
  wire                CsrAccessPlugin_logic_fsm_inject_trap;
  reg                 CsrAccessPlugin_logic_fsm_inject_unfreeze;
  wire                CsrAccessPlugin_logic_fsm_inject_freeze;
  reg                 CsrAccessPlugin_logic_fsm_inject_flushReg;
  wire                when_CsrAccessPlugin_l197;
  reg                 CsrAccessPlugin_logic_fsm_inject_sampled;
  reg                 CsrAccessPlugin_logic_fsm_inject_trapReg;
  reg                 CsrAccessPlugin_logic_fsm_inject_busTrapReg;
  reg        [3:0]    CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg;
  reg                 CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  reg                 CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo;
  wire                when_CsrAccessPlugin_l252;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  wire                when_CsrAccessPlugin_l279;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_mask;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_masked;
  wire       [31:0]   CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
  reg                 CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  reg                 CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo;
  wire                when_CsrAccessPlugin_l346;
  wire       [1:0]    switch_PrivilegedPlugin_l549;
  wire                when_CsrAccessPlugin_l346_1;
  wire                when_CsrAccessPlugin_l353;
  wire                when_CsrAccessPlugin_l346_2;
  wire                when_CsrAccessPlugin_l346_3;
  wire                when_CsrAccessPlugin_l346_4;
  wire                when_CsrAccessPlugin_l346_5;
  wire                when_CsrAccessPlugin_l346_6;
  wire                when_CsrAccessPlugin_l346_7;
  wire                when_CsrAccessPlugin_l346_8;
  wire                when_CsrAccessPlugin_l346_9;
  wire                when_CsrAccessPlugin_l346_10;
  wire                when_CsrAccessPlugin_l346_11;
  wire                when_CsrAccessPlugin_l343;
  wire                when_CsrAccessPlugin_l343_1;
  wire                when_CsrAccessPlugin_l346_12;
  wire                when_CsrAccessPlugin_l346_13;
  wire                when_CsrAccessPlugin_l346_14;
  wire                when_CsrAccessPlugin_l343_2;
  wire                when_CsrAccessPlugin_l343_3;
  wire                when_PerformanceCounterPlugin_l357;
  wire                when_PerformanceCounterPlugin_l359;
  wire       [31:0]   FetchL1Plugin_pmaBuilder_addressBits;
  wire                _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit;
  wire                FetchL1Plugin_pmaBuilder_onTransfers_0_hit;
  wire       [31:0]   LsuPlugin_pmaBuilder_l1_addressBits;
  wire       [0:0]    LsuPlugin_pmaBuilder_l1_argsBits;
  wire                _zz_LsuPlugin_logic_onPma_cached_rsp_io;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit;
  wire                LsuPlugin_pmaBuilder_l1_onTransfers_0_hit;
  wire       [31:0]   LsuPlugin_pmaBuilder_io_addressBits;
  wire       [2:0]    LsuPlugin_pmaBuilder_io_argsBits;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_0_hit;
  wire                _zz_LsuPlugin_logic_onPma_io_rsp_io;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_1_argsHit;
  wire                LsuPlugin_pmaBuilder_io_onTransfers_1_hit;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_hits;
  wire                CsrRamPlugin_logic_writeLogic_hit;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_input;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_oh;
  wire                CsrRamPlugin_logic_writeLogic_port_valid;
  wire       [3:0]    CsrRamPlugin_logic_writeLogic_port_payload_address;
  wire       [31:0]   CsrRamPlugin_logic_writeLogic_port_payload_data;
  wire                _zz_PerformanceCounterPlugin_logic_writePort_ready;
  wire                _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready;
  wire                _zz_CsrRamPlugin_csrMapper_write_ready;
  wire                _zz_CsrRamPlugin_setup_initPort_ready;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_hits;
  wire                CsrRamPlugin_logic_readLogic_hit;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_input;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  wire       [2:0]    CsrRamPlugin_logic_readLogic_oh;
  wire                _zz_CsrRamPlugin_logic_readLogic_sel;
  wire                _zz_CsrRamPlugin_logic_readLogic_sel_1;
  wire       [1:0]    CsrRamPlugin_logic_readLogic_sel;
  wire                CsrRamPlugin_logic_readLogic_port_cmd_valid;
  wire       [3:0]    CsrRamPlugin_logic_readLogic_port_cmd_payload;
  wire       [31:0]   CsrRamPlugin_logic_readLogic_port_rsp;
  reg        [2:0]    CsrRamPlugin_logic_readLogic_ohReg;
  reg                 CsrRamPlugin_logic_readLogic_busy;
  reg        [4:0]    CsrRamPlugin_logic_flush_counter;
  wire                CsrRamPlugin_logic_flush_done;
  wire                execute_lane0_bypasser_integer_RS1_port_valid;
  wire       [4:0]    execute_lane0_bypasser_integer_RS1_port_address;
  wire       [31:0]   execute_lane0_bypasser_integer_RS1_port_data;
  reg        [4:0]    execute_lane0_bypasser_integer_RS1_bypassEnables;
  wire       [4:0]    _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4;
  reg        [4:0]    _zz_execute_lane0_bypasser_integer_RS1_sel;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2;
  wire                execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3;
  wire       [4:0]    execute_lane0_bypasser_integer_RS1_sel;
  wire       [3:0]    _zz_execute_ctrl1_down_integer_RS1_lane0;
  (* keep , syn_keep *) reg        [31:0]   _zz_execute_ctrl1_down_integer_RS1_lane0_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l196;
  wire                execute_lane0_bypasser_integer_RS2_port_valid;
  wire       [4:0]    execute_lane0_bypasser_integer_RS2_port_address;
  wire       [31:0]   execute_lane0_bypasser_integer_RS2_port_data;
  reg        [4:0]    execute_lane0_bypasser_integer_RS2_bypassEnables;
  wire       [4:0]    _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4;
  reg        [4:0]    _zz_execute_lane0_bypasser_integer_RS2_sel;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2;
  wire                execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3;
  wire       [4:0]    execute_lane0_bypasser_integer_RS2_sel;
  wire       [3:0]    _zz_execute_ctrl1_down_integer_RS2_lane0;
  (* keep , syn_keep *) reg        [31:0]   _zz_execute_ctrl1_down_integer_RS2_lane0_1 /* synthesis syn_keep = 1 */ ;
  wire                when_ExecuteLanePlugin_l196_1;
  wire                execute_lane0_logic_completions_onCtrl_0_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_0_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_0_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_0_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_1_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_1_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_1_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_1_port_payload_commit;
  wire                execute_lane0_logic_completions_onCtrl_2_port_valid;
  wire       [15:0]   execute_lane0_logic_completions_onCtrl_2_port_payload_uopId;
  wire                execute_lane0_logic_completions_onCtrl_2_port_payload_trap;
  wire                execute_lane0_logic_completions_onCtrl_2_port_payload_commit;
  wire       [31:0]   execute_lane0_logic_decoding_decodingBits;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
  wire                _zz_execute_ctrl1_down_AguPlugin_SEL_lane0;
  wire                _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0;
  wire                _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1;
  wire                _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2;
  wire                _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
  wire                _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  wire                _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
  wire                _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  wire       [1:0]    _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  wire                _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2;
  wire                _zz_execute_ctrl1_down_AguPlugin_STORE_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1;
  wire       [1:0]    _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2;
  wire       [0:0]    _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0;
  wire       [0:0]    _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_1;
  wire       [0:0]    _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_2;
  wire                _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
  wire                _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
  wire       [2:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1;
  wire       [2:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  wire       [2:0]    _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3;
  wire                when_ExecuteLanePlugin_l306;
  wire                when_ExecuteLanePlugin_l306_1;
  wire                when_ExecuteLanePlugin_l306_2;
  wire                when_ExecuteLanePlugin_l306_3;
  wire                when_ExecuteLanePlugin_l306_4;
  wire                WhiteboxerPlugin_logic_csr_port_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_csr_port_payload_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_csr_port_payload_address;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_port_payload_write;
  wire       [31:0]   WhiteboxerPlugin_logic_csr_port_payload_read;
  wire                WhiteboxerPlugin_logic_csr_port_payload_writeDone;
  wire                WhiteboxerPlugin_logic_csr_port_payload_readDone;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_0_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_0_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_0_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_1_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_1_payload_data;
  wire                WhiteboxerPlugin_logic_rfWrites_ports_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_rfWrites_ports_2_payload_uopId;
  wire       [31:0]   WhiteboxerPlugin_logic_rfWrites_ports_2_payload_data;
  wire                WhiteboxerPlugin_logic_completions_ports_0_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_0_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_0_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_0_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_1_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_1_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_1_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_2_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_2_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_2_payload_commit;
  wire                WhiteboxerPlugin_logic_completions_ports_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_completions_ports_3_payload_uopId;
  wire                WhiteboxerPlugin_logic_completions_ports_3_payload_trap;
  wire                WhiteboxerPlugin_logic_completions_ports_3_payload_commit;
  wire                WhiteboxerPlugin_logic_commits_ports_0_oh_0;
  wire                WhiteboxerPlugin_logic_commits_ports_0_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_0_pc;
  wire       [31:0]   WhiteboxerPlugin_logic_commits_ports_0_uop;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_0_valid;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_0_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_1_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_1_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_1_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_2_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_2_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_2_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_3_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_3_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_3_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_4_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_4_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_4_payload_self;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_5_valid;
  wire       [15:0]   WhiteboxerPlugin_logic_reschedules_flushes_5_payload_uopId;
  wire                WhiteboxerPlugin_logic_reschedules_flushes_5_payload_self;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_valid;
  wire       [31:0]   early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice;
  wire       [31:0]   early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong;
  wire                early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget;
  wire       [11:0]   early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history;
  wire       [15:0]   early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId;
  wire       [1:0]    early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_valid;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_pcOnLastSlice;
  wire       [31:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_pcTarget;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_taken;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isBranch;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isPush;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_isPop;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_wasWrong;
  wire                WhiteboxerPlugin_logic_prediction_learns_0_payload_badPredictedTarget;
  wire       [11:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_history;
  wire       [15:0]   WhiteboxerPlugin_logic_prediction_learns_0_payload_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  wire                WhiteboxerPlugin_logic_loadExecute_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_loadExecute_uopId;
  wire       [1:0]    WhiteboxerPlugin_logic_loadExecute_size;
  wire       [31:0]   WhiteboxerPlugin_logic_loadExecute_address;
  wire       [31:0]   WhiteboxerPlugin_logic_loadExecute_data;
  wire                WhiteboxerPlugin_logic_storeCommit_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_storeCommit_uopId;
  wire       [11:0]   WhiteboxerPlugin_logic_storeCommit_storeId;
  wire       [1:0]    WhiteboxerPlugin_logic_storeCommit_size;
  wire       [31:0]   WhiteboxerPlugin_logic_storeCommit_address;
  wire       [31:0]   WhiteboxerPlugin_logic_storeCommit_data;
  wire                WhiteboxerPlugin_logic_storeCommit_amo;
  wire                WhiteboxerPlugin_logic_storeConditional_fire;
  wire       [15:0]   WhiteboxerPlugin_logic_storeConditional_uopId;
  wire                WhiteboxerPlugin_logic_storeConditional_miss;
  wire                WhiteboxerPlugin_logic_storeBroadcast_fire;
  wire       [11:0]   WhiteboxerPlugin_logic_storeBroadcast_storeId;
  wire                integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  wire       [4:0]    integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  wire       [31:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  wire       [15:0]   integer_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  reg        [5:0]    integer_RegFilePlugin_logic_initalizer_counter;
  wire                integer_RegFilePlugin_logic_initalizer_done;
  wire                when_RegFilePlugin_l130;
  wire                integer_write_0_valid /* verilator public */ ;
  wire       [4:0]    integer_write_0_address /* verilator public */ ;
  wire       [31:0]   integer_write_0_data /* verilator public */ ;
  wire       [15:0]   integer_write_0_uopId /* verilator public */ ;
  wire       [0:0]    WhiteboxerPlugin_logic_wfi;
  wire                WhiteboxerPlugin_logic_perf_executeFreezed;
  wire                WhiteboxerPlugin_logic_perf_dispatchHazards;
  wire       [0:0]    WhiteboxerPlugin_logic_perf_candidatesCount;
  wire       [0:0]    WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  reg                 _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  wire                when_Utils_l586;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  wire                when_Utils_l586_1;
  reg                 _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  wire                when_Utils_l586_2;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  wire                when_Utils_l586_3;
  reg                 _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
  reg        [59:0]   _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2;
  wire       [59:0]   WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  wire                WhiteboxerPlugin_logic_trap_ports_0_valid;
  wire                WhiteboxerPlugin_logic_trap_ports_0_interrupt;
  wire       [3:0]    WhiteboxerPlugin_logic_trap_ports_0_cause;
  wire                fetch_logic_ctrls_2_up_forgetOne;
  wire                fetch_logic_ctrls_1_up_forgetOne;
  wire                when_CtrlLink_l150;
  wire                when_CtrlLink_l157;
  wire                when_StageLink_l67;
  wire                when_DecodePipelinePlugin_l70;
  reg        [1:0]    LsuPlugin_logic_flusher_stateReg;
  reg        [1:0]    LsuPlugin_logic_flusher_stateNext;
  wire                when_LsuPlugin_l363;
  wire                when_LsuPlugin_l371;
  wire                LsuPlugin_logic_flusher_onExit_IDLE;
  wire                LsuPlugin_logic_flusher_onExit_CMD;
  wire                LsuPlugin_logic_flusher_onExit_COMPLETION;
  wire                LsuPlugin_logic_flusher_onEntry_IDLE;
  wire                LsuPlugin_logic_flusher_onEntry_CMD;
  wire                LsuPlugin_logic_flusher_onEntry_COMPLETION;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_stateReg;
  reg        [3:0]    TrapPlugin_logic_harts_0_trap_fsm_stateNext;
  wire                when_TrapPlugin_l409;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address;
  reg        [3:0]    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1;
  wire                when_TrapPlugin_l654;
  wire       [1:0]    switch_TrapPlugin_l655;
  wire                when_TrapPlugin_l509;
  wire       [2:0]    switch_TrapPlugin_l511;
  wire                when_TrapPlugin_l362;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_RESET;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_RUNNING;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_PROCESS_1;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVAL;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVEC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_ATS_RSP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_JUMP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_LSU_FLUSH;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onExit_FETCH_FLUSH;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_RESET;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_RUNNING;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_PROCESS_1;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVAL;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVEC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_EPC;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_APPLY;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_ATS_RSP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_JUMP;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_LSU_FLUSH;
  wire                TrapPlugin_logic_harts_0_trap_fsm_onEntry_FETCH_FLUSH;
  reg        [2:0]    MmuPlugin_logic_refill_stateReg;
  reg        [2:0]    MmuPlugin_logic_refill_stateNext;
  wire                when_MmuPlugin_l470;
  wire                when_MmuPlugin_l470_1;
  wire                when_MmuPlugin_l479;
  wire                when_MmuPlugin_l455;
  wire                _zz_57;
  wire                when_MmuPlugin_l455_1;
  wire                when_MmuPlugin_l487;
  wire                when_MmuPlugin_l455_2;
  wire                when_MmuPlugin_l455_3;
  wire                MmuPlugin_logic_refill_onExit_BOOT;
  wire                MmuPlugin_logic_refill_onExit_IDLE;
  wire                MmuPlugin_logic_refill_onExit_CMD_0;
  wire                MmuPlugin_logic_refill_onExit_CMD_1;
  wire                MmuPlugin_logic_refill_onExit_RSP_0;
  wire                MmuPlugin_logic_refill_onExit_RSP_1;
  wire                MmuPlugin_logic_refill_onEntry_BOOT;
  wire                MmuPlugin_logic_refill_onEntry_IDLE;
  wire                MmuPlugin_logic_refill_onEntry_CMD_0;
  wire                MmuPlugin_logic_refill_onEntry_CMD_1;
  wire                MmuPlugin_logic_refill_onEntry_RSP_0;
  wire                MmuPlugin_logic_refill_onEntry_RSP_1;
  reg        [2:0]    PerformanceCounterPlugin_logic_fsm_stateReg;
  reg        [2:0]    PerformanceCounterPlugin_logic_fsm_stateNext;
  wire                when_PerformanceCounterPlugin_l271;
  wire                when_PerformanceCounterPlugin_l278;
  wire                when_PerformanceCounterPlugin_l249;
  wire                when_PerformanceCounterPlugin_l255;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_BOOT;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_IDLE;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_READ_LOW;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_CALC_LOW;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_READ_HIGH;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_CALC_HIGH;
  wire                PerformanceCounterPlugin_logic_fsm_onExit_CSR_WRITE;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_BOOT;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_IDLE;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_READ_LOW;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_CALC_LOW;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_READ_HIGH;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_CALC_HIGH;
  wire                PerformanceCounterPlugin_logic_fsm_onEntry_CSR_WRITE;
  reg        [1:0]    CsrAccessPlugin_logic_fsm_stateReg;
  reg        [1:0]    CsrAccessPlugin_logic_fsm_stateNext;
  wire                when_CsrAccessPlugin_l296;
  wire                when_CsrAccessPlugin_l325;
  wire                when_CsrAccessPlugin_l212;
  wire                CsrAccessPlugin_logic_fsm_onExit_IDLE;
  wire                CsrAccessPlugin_logic_fsm_onExit_READ;
  wire                CsrAccessPlugin_logic_fsm_onExit_WRITE;
  wire                CsrAccessPlugin_logic_fsm_onExit_COMPLETION;
  wire                CsrAccessPlugin_logic_fsm_onEntry_IDLE;
  wire                CsrAccessPlugin_logic_fsm_onEntry_READ;
  wire                CsrAccessPlugin_logic_fsm_onEntry_WRITE;
  wire                CsrAccessPlugin_logic_fsm_onEntry_COMPLETION;
  `ifndef SYNTHESIS
  reg [31:0] execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [79:0] execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string;
  reg [39:0] execute_ctrl2_up_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string;
  reg [31:0] execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [79:0] execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string;
  reg [39:0] execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string;
  reg [31:0] execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [31:0] execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [39:0] execute_ctrl2_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string;
  reg [31:0] execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [79:0] execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string;
  reg [39:0] execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [127:0] FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string;
  reg [119:0] FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string;
  reg [95:0] LsuPlugin_logic_onAddress0_ls_port_payload_op_string;
  reg [95:0] LsuPlugin_logic_onAddress0_access_port_payload_op_string;
  reg [95:0] LsuPlugin_logic_onAddress0_flush_port_payload_op_string;
  reg [127:0] LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string;
  reg [119:0] LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string;
  reg [127:0] LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string;
  reg [119:0] LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string;
  reg [127:0] _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string;
  reg [39:0] _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string;
  reg [39:0] _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string;
  reg [39:0] _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string;
  reg [31:0] _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string;
  reg [39:0] _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string;
  reg [39:0] _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_1_string;
  reg [39:0] _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_2_string;
  reg [79:0] _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string;
  reg [79:0] _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string;
  reg [79:0] _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string;
  reg [79:0] LsuPlugin_logic_flusher_stateReg_string;
  reg [79:0] LsuPlugin_logic_flusher_stateNext_string;
  reg [87:0] TrapPlugin_logic_harts_0_trap_fsm_stateReg_string;
  reg [87:0] TrapPlugin_logic_harts_0_trap_fsm_stateNext_string;
  reg [39:0] MmuPlugin_logic_refill_stateReg_string;
  reg [39:0] MmuPlugin_logic_refill_stateNext_string;
  reg [71:0] PerformanceCounterPlugin_logic_fsm_stateReg_string;
  reg [71:0] PerformanceCounterPlugin_logic_fsm_stateNext_string;
  reg [79:0] CsrAccessPlugin_logic_fsm_stateReg_string;
  reg [79:0] CsrAccessPlugin_logic_fsm_stateNext_string;
  `endif

  reg [63:0] FetchL1Plugin_logic_banks_0_mem [0:511];
  reg [63:0] FetchL1Plugin_logic_banks_1_mem [0:511];
  reg [63:0] FetchL1Plugin_logic_banks_2_mem [0:511];
  reg [63:0] FetchL1Plugin_logic_banks_3_mem [0:511];
  reg [21:0] FetchL1Plugin_logic_ways_0_mem [0:63];
  reg [21:0] FetchL1Plugin_logic_ways_1_mem [0:63];
  reg [21:0] FetchL1Plugin_logic_ways_2_mem [0:63];
  reg [21:0] FetchL1Plugin_logic_ways_3_mem [0:63];
  reg [2:0] FetchL1Plugin_logic_plru_mem [0:63];
  reg [1:0] GSharePlugin_logic_mem_counter [0:16383];
  (* ram_style = "block" *) reg [48:0] BtbPlugin_logic_mem [0:511];
  reg [21:0] LsuL1Plugin_logic_ways_0_mem [0:63];
  reg [21:0] LsuL1Plugin_logic_ways_1_mem [0:63];
  reg [21:0] LsuL1Plugin_logic_ways_2_mem [0:63];
  reg [21:0] LsuL1Plugin_logic_ways_3_mem [0:63];
  reg [6:0] LsuL1Plugin_logic_shared_mem [0:63];
  reg [63:0] LsuL1Plugin_logic_writeback_victimBuffer [0:7];
  reg [31:0] CsrRamPlugin_logic_mem [0:15];
  function [2:0] zz_FetchL1Plugin_logic_trapPort_payload_arg(input dummy);
    begin
      zz_FetchL1Plugin_logic_trapPort_payload_arg = 3'b000;
      zz_FetchL1Plugin_logic_trapPort_payload_arg[1 : 0] = 2'b10;
      zz_FetchL1Plugin_logic_trapPort_payload_arg[2 : 2] = 1'b0;
    end
  endfunction
  wire [2:0] _zz_66;

  assign _zz_when = (! FetchL1Plugin_logic_refill_slots_0_valid);
  assign _zz_early0_IntAluPlugin_logic_alu_result = (early0_IntAluPlugin_logic_alu_bitwise | _zz_early0_IntAluPlugin_logic_alu_result_1);
  assign _zz_early0_IntAluPlugin_logic_alu_result_1 = (execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 ? execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 : 32'h0);
  assign _zz_early0_IntAluPlugin_logic_alu_result_2 = (execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0 ? _zz_early0_IntAluPlugin_logic_alu_result_3 : 32'h0);
  assign _zz_early0_IntAluPlugin_logic_alu_result_3 = _zz_early0_IntAluPlugin_logic_alu_result_4;
  assign _zz_early0_IntAluPlugin_logic_alu_result_5 = execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
  assign _zz_early0_IntAluPlugin_logic_alu_result_4 = {31'd0, _zz_early0_IntAluPlugin_logic_alu_result_5};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_amplitude = execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[4 : 0];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[0],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[1],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[2],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[3],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[4],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[5],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[6],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[7],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[8],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_1,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_2,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_3}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_shifted = ($signed(_zz_early0_BarrelShifterPlugin_logic_shift_shifted_1) >>> early0_BarrelShifterPlugin_logic_shift_amplitude);
  assign _zz_early0_BarrelShifterPlugin_logic_shift_shifted_1 = {(execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0 && execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]),early0_BarrelShifterPlugin_logic_shift_reversed};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched = {early0_BarrelShifterPlugin_logic_shift_shifted[0],{early0_BarrelShifterPlugin_logic_shift_shifted[1],{early0_BarrelShifterPlugin_logic_shift_shifted[2],{early0_BarrelShifterPlugin_logic_shift_shifted[3],{early0_BarrelShifterPlugin_logic_shift_shifted[4],{early0_BarrelShifterPlugin_logic_shift_shifted[5],{early0_BarrelShifterPlugin_logic_shift_shifted[6],{early0_BarrelShifterPlugin_logic_shift_shifted[7],{early0_BarrelShifterPlugin_logic_shift_shifted[8],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_1,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_2,_zz_early0_BarrelShifterPlugin_logic_shift_patched_3}}}}}}}}}}};
  assign _zz_execute_ctrl2_down_MUL_SRC1_lane0 = {(execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 && execute_ctrl2_up_integer_RS1_lane0[31]),execute_ctrl2_up_integer_RS1_lane0};
  assign _zz_execute_ctrl2_down_MUL_SRC2_lane0 = {(execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 && execute_ctrl2_up_integer_RS2_lane0[31]),execute_ctrl2_up_integer_RS2_lane0};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = {{13{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_1[33]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_2 = {1'b0,execute_ctrl2_down_MUL_SRC1_lane0[16 : 0]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0_3 = execute_ctrl2_down_MUL_SRC2_lane0[32 : 17];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = {{13{_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_1[33]}}, _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_1};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_2 = execute_ctrl2_down_MUL_SRC1_lane0[32 : 17];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0_3 = {1'b0,execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]};
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_1 = ($signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_2) * $signed(_zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_3));
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_1[29:0];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_2 = execute_ctrl2_down_MUL_SRC1_lane0[32 : 17];
  assign _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0_3 = execute_ctrl2_down_MUL_SRC2_lane0[32 : 17];
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_4 = {2'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_5 = {2'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6 = {2'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5);
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_4 = {2'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_5 = {2'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1};
  assign _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6 = {2'd0, _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2};
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1 = execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0;
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0 = {31'd0, _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0_1};
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1 = execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0;
  assign _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0 = {31'd0, _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0_1};
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1 = ((early0_DivPlugin_logic_processing_divRevertResult ? (~ _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0) : _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0) + _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2);
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3 = early0_DivPlugin_logic_processing_divRevertResult;
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_2 = {31'd0, _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_3};
  assign _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits = (fetch_logic_ctrls_1_down_Fetch_WORD_PC >>> 4'd12);
  assign _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits = (fetch_logic_ctrls_1_down_Fetch_WORD_PC >>> 4'd12);
  assign _zz_FetchL1Plugin_logic_hits_w_2_indirect_bypassHits = (fetch_logic_ctrls_1_down_Fetch_WORD_PC >>> 4'd12);
  assign _zz_FetchL1Plugin_logic_hits_w_3_indirect_bypassHits = (fetch_logic_ctrls_1_down_Fetch_WORD_PC >>> 4'd12);
  assign _zz_FetchL1Plugin_logic_ctrl_dataAccessFault = (((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error : 1'b0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error : 1'b0)) | ((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_2 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_2_error : 1'b0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_3 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_3_error : 1'b0)));
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_5 = fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_4 = {2'd0, _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_5};
  assign _zz_BtbPlugin_logic_ras_ptr_push = (BtbPlugin_logic_ras_ptr_push + _zz_BtbPlugin_logic_ras_ptr_push_1);
  assign _zz_BtbPlugin_logic_ras_ptr_push_2 = BtbPlugin_logic_ras_ptr_pushIt;
  assign _zz_BtbPlugin_logic_ras_ptr_push_1 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_push_2};
  assign _zz_BtbPlugin_logic_ras_ptr_push_4 = BtbPlugin_logic_ras_ptr_popIt;
  assign _zz_BtbPlugin_logic_ras_ptr_push_3 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_push_4};
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue = (BtbPlugin_logic_ras_ptr_pop + _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1);
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2 = BtbPlugin_logic_ras_ptr_pushIt;
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_1 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_2};
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4 = BtbPlugin_logic_ras_ptr_popIt;
  assign _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3 = {1'd0, _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_4};
  assign _zz_WhiteboxerPlugin_logic_decodes_0_pc = {32'd0, decode_ctrls_0_down_PC_0};
  assign _zz_PerformanceCounterPlugin_logic_eventInstructions_0 = ((! PerformanceCounterPlugin_logic_ignoreNextCommit) ? PerformanceCounterPlugin_logic_commitMask : 1'b0);
  assign _zz_PerformanceCounterPlugin_logic_counters_cycle_value_1 = (! PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit);
  assign _zz_PerformanceCounterPlugin_logic_counters_cycle_value = {7'd0, _zz_PerformanceCounterPlugin_logic_counters_cycle_value_1};
  assign _zz_PerformanceCounterPlugin_logic_counters_instret_value_1 = {7'd0, _zz_PerformanceCounterPlugin_logic_counters_instret_value};
  assign _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl1_down_Decode_UOP_lane0[31 : 20];
  assign _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1 = {execute_ctrl1_down_Decode_UOP_lane0[31 : 25],execute_ctrl1_down_Decode_UOP_lane0[11 : 7]};
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 = ($signed(execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0) + $signed(early0_SrcPlugin_logic_addsub_combined_rs2Patched));
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1 = _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2;
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3 = execute_ctrl2_down_SrcStageables_REVERT_lane0;
  assign _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_2 = {31'd0, _zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_3};
  assign _zz_early0_BranchPlugin_pcCalc_target_b = {{{{execute_ctrl2_down_Decode_UOP_lane0[31],execute_ctrl2_down_Decode_UOP_lane0[19 : 12]},execute_ctrl2_down_Decode_UOP_lane0[20]},execute_ctrl2_down_Decode_UOP_lane0[30 : 21]},1'b0};
  assign _zz_early0_BranchPlugin_pcCalc_target_b_1 = execute_ctrl2_down_Decode_UOP_lane0[31 : 20];
  assign _zz_early0_BranchPlugin_pcCalc_target_b_2 = {{{{execute_ctrl2_down_Decode_UOP_lane0[31],execute_ctrl2_down_Decode_UOP_lane0[7]},execute_ctrl2_down_Decode_UOP_lane0[30 : 25]},execute_ctrl2_down_Decode_UOP_lane0[11 : 8]},1'b0};
  assign _zz_early0_BranchPlugin_pcCalc_slices_1 = 1'b0;
  assign _zz_early0_BranchPlugin_pcCalc_slices = {1'd0, _zz_early0_BranchPlugin_pcCalc_slices_1};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = ($signed(early0_BranchPlugin_pcCalc_target_a) + $signed(early0_BranchPlugin_pcCalc_target_b));
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1 = ({2'd0,early0_BranchPlugin_pcCalc_slices} <<< 2'd2);
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = {28'd0, _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0_1};
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1 = 2'b00;
  assign _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = {30'd0, _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0_1};
  assign _zz__zz_CfuPlugin_logic_bus_cmd_payload_inputs_1_1 = execute_ctrl2_down_Decode_UOP_lane0[31 : 24];
  assign _zz__zz_CfuPlugin_logic_bus_cmd_payload_inputs_1 = {{24{_zz__zz_CfuPlugin_logic_bus_cmd_payload_inputs_1_1[7]}}, _zz__zz_CfuPlugin_logic_bus_cmd_payload_inputs_1_1};
  assign _zz_early0_EnvPlugin_logic_trapPort_payload_code = {2'd0, early0_EnvPlugin_logic_exe_privilege};
  assign _zz_early0_BranchPlugin_logic_alu_expectedMsb = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
  assign _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_1 = {early0_BranchPlugin_logic_jumpLogic_history_shifter,execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0};
  assign _zz_decode_ctrls_1_down_RS1_ENABLE_0 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000044) == 32'h0),{_zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0,{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00006004) == 32'h00002000),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00005004) == 32'h00001000),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002050) == 32'h00002000)}}}});
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000002c) == 32'h00000008),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000054) == 32'h00000040),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000006c) == 32'h00000020),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RS2_ENABLE_0_1) == 32'h08002004),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RS2_ENABLE_0_2) == 32'h00002004)}}}});
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000048) == 32'h00000048),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001010) == 32'h00001010),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002010) == 32'h00002010),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_RD_ENABLE_0_1) == 32'h00002008),{(_zz_decode_ctrls_1_down_RD_ENABLE_0_2 == _zz_decode_ctrls_1_down_RD_ENABLE_0_3),{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0,{_zz_decode_ctrls_1_down_RD_ENABLE_0_4,_zz_decode_ctrls_1_down_RD_ENABLE_0_5}}}}}}});
  assign _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb = (|((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000050) == 32'h00000040));
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1 = ((! decode_ctrls_1_down_Prediction_ALIGN_REDO_0) ? 2'b00 : 2'b00);
  assign _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = {30'd0, _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice_1};
  assign _zz_GSharePlugin_logic_onLearn_hash_5 = LearnPlugin_logic_learn_payload_history;
  assign _zz_GSharePlugin_logic_onLearn_hash_4 = {2'd0, _zz_GSharePlugin_logic_onLearn_hash_5};
  assign _zz_BtbPlugin_logic_memWrite_payload_address = (LearnPlugin_logic_learn_payload_pcOnLastSlice >>> 2'd2);
  assign _zz_decode_ctrls_1_down_CfuPlugin_logic_CFU_ENABLE_0 = _zz_decode_ctrls_1_down_CfuPlugin_logic_CFU_ENABLE_0_1[0];
  assign _zz_decode_ctrls_1_down_CfuPlugin_logic_CFU_ENABLE_0_1 = (|_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0);
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1[0];
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0_1 = 1'b0;
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1[0];
  assign _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0_1 = 1'b0;
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_2[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_2 = (|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000040) == 32'h00000040),{_zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0,{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001014) == 32'h00001004),((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002014) == 32'h00002004)}}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0,{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0,{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0 = _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1});
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0_1 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0,{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1}});
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_4[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_4 = (|{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0,{_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2,_zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1}});
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0_1 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_2[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_2 = (|_zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0);
  assign _zz_BtbPlugin_logic_memWrite_payload_address_1 = (DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice >>> 2'd2);
  assign _zz_BtbPlugin_logic_memRead_cmd_payload = (fetch_logic_ctrls_0_down_Fetch_WORD_PC >>> 2'd2);
  assign _zz_BtbPlugin_logic_ras_write_payload_data = (BtbPlugin_logic_applyIt_rasLogic_pushPc + 32'h00000004);
  assign _zz_LsuL1Plugin_logic_writeback_read_wordIndex_1 = LsuL1Plugin_logic_writeback_read_slotRead_valid;
  assign _zz_LsuL1Plugin_logic_writeback_read_wordIndex = {2'd0, _zz_LsuL1Plugin_logic_writeback_read_wordIndex_1};
  assign _zz_LsuL1Plugin_logic_writeback_write_wordIndex_1 = (LsuL1Plugin_logic_writeback_write_bufferRead_fire && 1'b1);
  assign _zz_LsuL1Plugin_logic_writeback_write_wordIndex = {2'd0, _zz_LsuL1Plugin_logic_writeback_write_wordIndex_1};
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback = ({execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded,{execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded,{execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded,execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded}}} & execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty);
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_doWrite = (((_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 ? (1'b1 && (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault)) : 1'b0) | (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 ? (1'b1 && (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault)) : 1'b0)) | ((_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_2 ? (1'b1 && (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault)) : 1'b0) | (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_3 ? (1'b1 && (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault)) : 1'b0)));
  assign _zz_58 = (_zz_59 + _zz_61);
  assign _zz_63 = _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_3;
  assign _zz_62 = {2'd0, _zz_63};
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty_1 = (4'b0001 <<< LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate);
  assign _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1 = ({2'd0,TrapPlugin_logic_harts_0_trap_fsm_jumpOffset} <<< 2'd2);
  assign _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget = {29'd0, _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget_1};
  assign _zz_LsuPlugin_logic_onAddress0_ls_storeId_1 = LsuPlugin_logic_onAddress0_ls_port_fire;
  assign _zz_LsuPlugin_logic_onAddress0_ls_storeId = {11'd0, _zz_LsuPlugin_logic_onAddress0_ls_storeId_1};
  assign _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address = ({6'd0,LsuPlugin_logic_flusher_cmdCounter} <<< 3'd6);
  assign _zz_LsuPlugin_logic_onPma_addressExtension = execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub = ($signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1) + $signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4));
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_1 = ($signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2) + $signed(_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3));
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_2 = execute_ctrl4_down_integer_RS2_lane0;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_3 = (LsuPlugin_logic_onCtrl_rva_alu_compare ? (~ LsuPlugin_logic_onCtrl_rva_srcBuffer) : LsuPlugin_logic_onCtrl_rva_srcBuffer);
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5 = (LsuPlugin_logic_onCtrl_rva_alu_compare ? 2'b01 : 2'b00);
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_4 = {{30{_zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5[1]}}, _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub_5};
  assign _zz_LsuPlugin_logic_onCtrl_rva_lrsc_age_1 = (! execute_freeze_valid);
  assign _zz_LsuPlugin_logic_onCtrl_rva_lrsc_age = {5'd0, _zz_LsuPlugin_logic_onCtrl_rva_lrsc_age_1};
  assign _zz_LsuPlugin_logic_trapPort_payload_code = (execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 ? (execute_ctrl4_down_LsuL1_STORE_lane0 ? 3'b110 : 3'b100) : 3'b000);
  assign _zz_LsuPlugin_logic_flusher_cmdCounter = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign _zz_PcPlugin_logic_harts_0_self_pc_1 = (PcPlugin_logic_harts_0_self_increment ? 3'b100 : 3'b000);
  assign _zz_PcPlugin_logic_harts_0_self_pc = {29'd0, _zz_PcPlugin_logic_harts_0_self_pc_1};
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault = (((_zz_PcPlugin_logic_harts_0_aggregator_target ? TrapPlugin_logic_harts_0_trap_pcPort_payload_fault : 1'b0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_1 ? early0_BranchPlugin_logic_pcPort_payload_fault : 1'b0)) | (_zz_PcPlugin_logic_harts_0_aggregator_target_2 ? PcPlugin_logic_harts_0_self_flow_payload_fault : 1'b0));
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault_1_1 = (_zz_PcPlugin_logic_harts_0_aggregator_fault_1 ? BtbPlugin_logic_pcPort_payload_fault : 1'b0);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext_1 = LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement;
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = {1'd0, _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext_1};
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_4 = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowExecute : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowExecute : 1'b0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowExecute : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowExecute : 1'b0)));
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowRead : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowRead : 1'b0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowRead : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowRead : 1'b0)));
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowWrite : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowWrite : 1'b0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowWrite : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowWrite : 1'b0)));
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowUser : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowUser : 1'b0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowUser : 1'b0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowUser : 1'b0)));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_3 = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowExecute : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowExecute : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowExecute : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowRead : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowRead : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowRead : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowWrite : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowWrite : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowWrite : 1'b0));
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowUser : 1'b0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowUser : 1'b0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowUser : 1'b0));
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_a = PerformanceCounterPlugin_logic_fsm_counterReaded[6:0];
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_b = ({7'd0,PerformanceCounterPlugin_logic_fsm_counterReaded[7]} <<< 3'd7);
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_sum_1 = {1'b0,PerformanceCounterPlugin_logic_fsm_calc_b};
  assign _zz_PerformanceCounterPlugin_logic_fsm_calc_sum = {24'd0, _zz_PerformanceCounterPlugin_logic_fsm_calc_sum_1};
  assign _zz_PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked = (PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input - 2'b01);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23 = ({19'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue ? MmuPlugin_logic_status_mxr : 1'b0)} <<< 5'd19);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22 = {12'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_23};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25 = ({18'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue ? MmuPlugin_logic_status_sum : 1'b0)} <<< 5'd18);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24 = {13'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_25};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28 = ({19'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? MmuPlugin_logic_status_mxr : 1'b0)} <<< 5'd19);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 = {12'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_28};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30 = ({18'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 ? MmuPlugin_logic_status_sum : 1'b0)} <<< 5'd18);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29 = {13'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_30};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 ? MmuPlugin_logic_satp_mode : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 ? MmuPlugin_logic_satp_ppn : 20'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34 = {12'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_35};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? CfuPlugin_logic_en : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39 = ({16'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? CfuPlugin_logic_csr_stateId : 3'b000)} <<< 5'd16);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38 = {13'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_39};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 ? CfuPlugin_logic_csr_cfuIndex : 4'b0000);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_43};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46 = ((when_CsrService_l198 && REG_CSR_3858) ? 6'h2e : 6'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_46};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_status_mpie : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_51};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_status_mie : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_53};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_57 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_status_mpp : 2'b00)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56 = {19'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_57};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_58 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_status_sd : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_61 = ({17'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_status_mprv : 1'b0)} <<< 5'd17);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_60 = {14'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_61};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_63 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_status_fs : 2'b00)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_62 = {17'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_63};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_67 = ({22'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_status_tsr : 1'b0)} <<< 5'd22);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_66 = {9'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_67};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_69 = ({20'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_status_tvm : 1'b0)} <<< 5'd20);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_68 = {11'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_69};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_72 = ({21'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_m_status_tw : 1'b0)} <<< 5'd21);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_71 = {10'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_72};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_73 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PrivilegedPlugin_logic_harts_0_m_cause_interrupt : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_77 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 ? PrivilegedPlugin_logic_harts_0_m_cause_code : 4'b0000);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_76 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_77};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_79 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 ? PrivilegedPlugin_logic_harts_0_m_ip_meip : 1'b0)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_78 = {20'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_79};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_82 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 ? PrivilegedPlugin_logic_harts_0_m_ip_mtip : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_81 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_82};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_84 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 ? PrivilegedPlugin_logic_harts_0_m_ip_msip : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_83 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_84};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_88 = ({11'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_m_ie_meie : 1'b0)} <<< 4'd11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_87 = {20'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_88};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_90 = ({7'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_m_ie_mtie : 1'b0)} <<< 3'd7);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_89 = {24'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_90};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_93 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_m_ie_msie : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_92 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_93};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_95 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? PrivilegedPlugin_logic_harts_0_m_edeleg_iam : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_94 = {31'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_95};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_99 = ({3'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? PrivilegedPlugin_logic_harts_0_m_edeleg_bp : 1'b0)} <<< 2'd3);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_98 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_99};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_101 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? PrivilegedPlugin_logic_harts_0_m_edeleg_eu : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_100 = {23'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_101};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_104 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? PrivilegedPlugin_logic_harts_0_m_edeleg_es : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_103 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_104};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_106 = ({12'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? PrivilegedPlugin_logic_harts_0_m_edeleg_ipf : 1'b0)} <<< 4'd12);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_105 = {19'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_106};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_110 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? PrivilegedPlugin_logic_harts_0_m_edeleg_lpf : 1'b0)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_109 = {18'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_110};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_112 = ({15'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 ? PrivilegedPlugin_logic_harts_0_m_edeleg_spf : 1'b0)} <<< 4'd15);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_111 = {16'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_112};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_115 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_ideleg_se : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_114 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_115};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_117 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_ideleg_st : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_116 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_117};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_121 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 ? PrivilegedPlugin_logic_harts_0_m_ideleg_ss : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_120 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_121};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_122 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 ? PrivilegedPlugin_logic_harts_0_s_cause_interrupt : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_125 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 ? PrivilegedPlugin_logic_harts_0_s_cause_code : 4'b0000);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_124 = {28'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_125};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_126 = ({31'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 ? PrivilegedPlugin_logic_harts_0_m_status_sd : 1'b0)} <<< 5'd31);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_130 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_s_status_spp : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_129 = {23'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_130};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_132 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_s_status_spie : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_131 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_132};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_135 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 ? PrivilegedPlugin_logic_harts_0_s_status_sie : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_134 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_135};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_137 = ({8'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 ? PrivilegedPlugin_logic_harts_0_s_status_spp : 1'b0)} <<< 4'd8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_136 = {23'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_137};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_141 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 ? PrivilegedPlugin_logic_harts_0_s_status_spie : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_140 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_141};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_143 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 ? PrivilegedPlugin_logic_harts_0_s_status_sie : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_142 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_143};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_146 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 ? PrivilegedPlugin_logic_harts_0_m_status_fs : 2'b00)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_145 = {17'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_146};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_148 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_s_ie_seie : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_147 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_148};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_152 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 ? (PrivilegedPlugin_logic_harts_0_s_ie_seie && PrivilegedPlugin_logic_harts_0_m_ideleg_se) : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_151 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_152};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_154 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_s_ie_stie : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_153 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_154};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_157 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 ? (PrivilegedPlugin_logic_harts_0_s_ie_stie && PrivilegedPlugin_logic_harts_0_m_ideleg_st) : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_156 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_157};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_159 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 ? PrivilegedPlugin_logic_harts_0_s_ie_ssie : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_158 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_159};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_163 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 ? (PrivilegedPlugin_logic_harts_0_s_ie_ssie && PrivilegedPlugin_logic_harts_0_m_ideleg_ss) : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_162 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_163};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_165 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 ? PrivilegedPlugin_logic_harts_0_s_ip_seipOr : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_164 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_165};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_168 = ({9'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 ? (PrivilegedPlugin_logic_harts_0_s_ip_seipOr && PrivilegedPlugin_logic_harts_0_m_ideleg_se) : 1'b0)} <<< 4'd9);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_167 = {22'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_168};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_170 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 ? PrivilegedPlugin_logic_harts_0_s_ip_stip : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_169 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_170};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_174 = ({5'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 ? (PrivilegedPlugin_logic_harts_0_s_ip_stip && PrivilegedPlugin_logic_harts_0_m_ideleg_st) : 1'b0)} <<< 3'd5);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_173 = {26'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_174};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_176 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 ? PrivilegedPlugin_logic_harts_0_s_ip_ssip : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_175 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_176};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_179 = ({1'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 ? (PrivilegedPlugin_logic_harts_0_s_ip_ssip && PrivilegedPlugin_logic_harts_0_m_ideleg_ss) : 1'b0)} <<< 1'd1);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_178 = {30'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_179};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_185 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 ? PerformanceCounterPlugin_logic_counters_cycle_mcounteren : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_184 = {31'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_185};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_187 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 ? PerformanceCounterPlugin_logic_counters_cycle_scounteren : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_186 = {31'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_187};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_189 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 ? PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit : 1'b0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_188 = {31'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_189};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_191 = ({2'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 ? PerformanceCounterPlugin_logic_counters_instret_mcounteren : 1'b0)} <<< 2'd2);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_190 = {29'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_191};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_193 = ({2'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 ? PerformanceCounterPlugin_logic_counters_instret_scounteren : 1'b0)} <<< 2'd2);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_192 = {29'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_193};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_195 = ({2'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 ? PerformanceCounterPlugin_logic_counters_instret_mcountinhibit : 1'b0)} <<< 2'd2);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_194 = {29'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_195};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_199 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 ? PerformanceCounterPlugin_logic_interrupt_ip : 1'b0)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_198 = {18'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_199};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_201 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 ? PerformanceCounterPlugin_logic_interrupt_ie : 1'b0)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_200 = {18'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_201};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_203 = ({13'd0,(_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 ? PerformanceCounterPlugin_logic_interrupt_sup_deleg : 1'b0)} <<< 4'd13);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_202 = {18'd0, _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_203};
  assign _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1 = CsrAccessPlugin_logic_fsm_interface_uop[19 : 15];
  assign _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = {27'd0, _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask_1};
  assign _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit = (|_zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io);
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io_1 = (|_zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io);
  assign _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit = (|_zz_LsuPlugin_logic_onPma_cached_rsp_io);
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_io_1 = (|_zz_LsuPlugin_logic_onPma_cached_rsp_io);
  assign _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit = (|{((LsuPlugin_pmaBuilder_io_addressBits & 32'h01800000) == 32'h00800000),((LsuPlugin_pmaBuilder_io_addressBits & 32'h01010000) == 32'h00010000)});
  assign _zz_LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit = (|{_zz_LsuPlugin_logic_onPma_io_rsp_io,((LsuPlugin_pmaBuilder_io_addressBits & 32'h00810000) == 32'h0)});
  assign _zz_LsuPlugin_logic_onPma_io_rsp_io_1 = (|_zz_LsuPlugin_logic_onPma_io_rsp_io);
  assign _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input - 4'b0001);
  assign _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input - 3'b001);
  assign _zz_CsrRamPlugin_logic_flush_counter_1 = (! CsrRamPlugin_logic_flush_done);
  assign _zz_CsrRamPlugin_logic_flush_counter = {4'd0, _zz_CsrRamPlugin_logic_flush_counter_1};
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00002030) == 32'h00002010),{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0,{((execute_lane0_logic_decoding_decodingBits & 32'h00001030) == 32'h00000010),{((execute_lane0_logic_decoding_decodingBits & 32'h02002050) == 32'h00002010),((execute_lane0_logic_decoding_decodingBits & 32'h02001050) == 32'h00000010)}}}});
  assign _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00003034) == 32'h00001010),((execute_lane0_logic_decoding_decodingBits & 32'h02003054) == 32'h00001010)});
  assign _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0_1 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0);
  assign _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h02004074) == 32'h02000030));
  assign _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h0200406c) == 32'h02004020));
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00001054) == 32'h00001004),((execute_lane0_logic_decoding_decodingBits & 32'h00003050) == 32'h00000050)});
  assign _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0 = _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0_1[0];
  assign _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0_1 = (|_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00001050) == 32'h00001050),((execute_lane0_logic_decoding_decodingBits & 32'h00002050) == 32'h00002050)});
  assign _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_1 = _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_2[0];
  assign _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_2 = (|{_zz_execute_ctrl1_down_AguPlugin_SEL_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h00001054) == 32'h00000004)});
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1[0];
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00003054) == 32'h00000004));
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1 = _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_2[0];
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00000048) == 32'h00000048),{((execute_lane0_logic_decoding_decodingBits & 32'h00001010) == 32'h00001010),{((execute_lane0_logic_decoding_decodingBits & 32'h00002010) == 32'h00002010),{_zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0,{(_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_3 == _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_4),{_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0,{_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_5,_zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_6}}}}}}});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1}}}}});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1}}});
  assign _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0_1[0];
  assign _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0}});
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_6 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1}}}}});
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_5 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1}}});
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_4[0];
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_4 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1,_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0}});
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_2[0];
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_2 = (|{_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0,_zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0});
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1[0];
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00006004) == 32'h00002000));
  assign _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0 = _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2,{((execute_lane0_logic_decoding_decodingBits & 32'h00002014) == 32'h00002010),((execute_lane0_logic_decoding_decodingBits & 32'h40000034) == 32'h40000030)}});
  assign _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0 = _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00000024) == 32'h00000024));
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00004010) == 32'h0));
  assign _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0_1[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0_1 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0,{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h02000068) == 32'h00000020)}}});
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_3 = _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_4[0];
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_4 = (|{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2,{((execute_lane0_logic_decoding_decodingBits & 32'h00004010) == 32'h00004010),{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1,{_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h02000028) == 32'h00000020)}}}});
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1[0];
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0_1 = (|{_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0,{((execute_lane0_logic_decoding_decodingBits & 32'h00000018) == 32'h0),((execute_lane0_logic_decoding_decodingBits & 32'h00002014) == 32'h00002004)}});
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1[0];
  assign _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0_1 = (|{_zz_execute_ctrl1_down_AguPlugin_SEL_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h00002054) == 32'h00002004)});
  assign _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0 = _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00002010) == 32'h00002000),((execute_lane0_logic_decoding_decodingBits & 32'h00005000) == 32'h00001000)});
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1 = _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_2 = (|_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0);
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h40000000) == 32'h40000000));
  assign _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0 = _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0_1[0];
  assign _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0_1 = (|{_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0,_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0});
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1[0];
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0_1 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00001000) == 32'h0),_zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0});
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_2[0];
  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h00005000) == 32'h00004000),_zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0});
  assign _zz_execute_ctrl1_down_DivPlugin_REM_lane0 = _zz_execute_ctrl1_down_DivPlugin_REM_lane0_1[0];
  assign _zz_execute_ctrl1_down_DivPlugin_REM_lane0_1 = (|_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00004000) == 32'h00004000));
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_2[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_2 = (|_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_2[0];
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_2 = (|_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0);
  assign _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_1 = _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_2[0];
  assign _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_2 = (|{_zz_execute_ctrl1_down_AguPlugin_LOAD_lane0,{((execute_lane0_logic_decoding_decodingBits & 32'h08002008) == 32'h00002008),((execute_lane0_logic_decoding_decodingBits & 32'h10002008) == 32'h00002008)}});
  assign _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_1 = _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_2[0];
  assign _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_2 = (|{((execute_lane0_logic_decoding_decodingBits & 32'h08000020) == 32'h08000020),{_zz_execute_ctrl1_down_AguPlugin_STORE_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h00000028) == 32'h00000020)}});
  assign _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1 = _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_2[0];
  assign _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_2 = (|_zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0);
  assign _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0 = _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0_1 = 1'b0;
  assign _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0 = _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0_1 = 1'b0;
  assign _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0 = _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0_1[0];
  assign _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0_1 = 1'b0;
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1[0];
  assign _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0_1 = 1'b0;
  assign _zz_WhiteboxerPlugin_logic_csr_access_payload_address = CsrAccessPlugin_logic_fsm_interface_uop;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1 = _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1_1};
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1;
  assign _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = {59'd0, _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1_1};
  assign _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = (2'b01 <<< FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = (MmuPlugin_logic_refill_storageOhReg[1] ? _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask_1 : 4'b0000);
  assign _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask_1 = (4'b0001 <<< LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value);
  assign _zz_PerformanceCounterPlugin_logic_writePort_data = PerformanceCounterPlugin_logic_fsm_calc_sum;
  assign _zz_PerformanceCounterPlugin_logic_writePort_data_1 = PerformanceCounterPlugin_logic_fsm_calc_sum;
  assign _zz_PerformanceCounterPlugin_logic_counters_cycle_value_2 = CsrAccessPlugin_bus_write_bits;
  assign _zz_PerformanceCounterPlugin_logic_counters_instret_value_2 = CsrAccessPlugin_bus_write_bits;
  assign _zz_FetchL1Plugin_logic_ways_0_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_0_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[0];
  assign _zz_FetchL1Plugin_logic_ways_1_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_1_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[1];
  assign _zz_FetchL1Plugin_logic_ways_2_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_2_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[2];
  assign _zz_FetchL1Plugin_logic_ways_3_mem_port = {FetchL1Plugin_logic_waysWrite_tag_address,{FetchL1Plugin_logic_waysWrite_tag_error,FetchL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_FetchL1Plugin_logic_ways_3_mem_port_1 = FetchL1Plugin_logic_waysWrite_mask[3];
  assign _zz_FetchL1Plugin_logic_plru_mem_port = {FetchL1Plugin_logic_plru_write_payload_data_1,FetchL1Plugin_logic_plru_write_payload_data_0};
  assign _zz_GSharePlugin_logic_mem_counter_port = GSharePlugin_logic_mem_write_payload_data_0;
  assign _zz_BtbPlugin_logic_mem_port = {BtbPlugin_logic_memDp_wp_payload_data_0_isPop,{BtbPlugin_logic_memDp_wp_payload_data_0_isPush,{BtbPlugin_logic_memDp_wp_payload_data_0_isBranch,{BtbPlugin_logic_memDp_wp_payload_data_0_pcTarget,BtbPlugin_logic_memDp_wp_payload_data_0_hash}}}};
  assign _zz_LsuL1Plugin_logic_ways_0_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_0_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[0];
  assign _zz_LsuL1Plugin_logic_ways_1_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_1_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[1];
  assign _zz_LsuL1Plugin_logic_ways_2_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_2_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[2];
  assign _zz_LsuL1Plugin_logic_ways_3_mem_port = {LsuL1Plugin_logic_waysWrite_tag_fault,{LsuL1Plugin_logic_waysWrite_tag_address,LsuL1Plugin_logic_waysWrite_tag_loaded}};
  assign _zz_LsuL1Plugin_logic_ways_3_mem_port_1 = LsuL1Plugin_logic_waysWrite_mask[3];
  assign _zz_LsuL1Plugin_logic_shared_mem_port = {LsuL1Plugin_logic_shared_write_payload_data_dirty,{LsuL1Plugin_logic_shared_write_payload_data_plru_1,LsuL1Plugin_logic_shared_write_payload_data_plru_0}};
  assign _zz_LsuL1Plugin_logic_writeback_victimBuffer_port = LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex;
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 2];
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 2];
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 2];
  assign _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[2 : 2];
  assign _zz_PerformanceCounterPlugin_logic_commitCount_1 = PerformanceCounterPlugin_logic_commitMask[0];
  assign _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0_1 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1_1 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2_1 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3_1 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[2 : 2];
  assign _zz_60 = {_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_2,{_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1,_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0}};
  assign _zz_65 = {_zz_53[2],{_zz_53[1],_zz_53[0]}};
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_1 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[1 : 0];
  assign _zz_LsuPlugin_logic_onCtrl_loadData_shifted_3 = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[1 : 1];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_0_2 = _zz_PerformanceCounterPlugin_logic_events_sums_0[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_1_2 = _zz_PerformanceCounterPlugin_logic_events_sums_1[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_2_2 = _zz_PerformanceCounterPlugin_logic_events_sums_2[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_3_2 = _zz_PerformanceCounterPlugin_logic_events_sums_3[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_4_2 = _zz_PerformanceCounterPlugin_logic_events_sums_4[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_5_2 = _zz_PerformanceCounterPlugin_logic_events_sums_5[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_6_2 = _zz_PerformanceCounterPlugin_logic_events_sums_6[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_7_2 = _zz_PerformanceCounterPlugin_logic_events_sums_7[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_8_2 = _zz_PerformanceCounterPlugin_logic_events_sums_8[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_9_2 = _zz_PerformanceCounterPlugin_logic_events_sums_9[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_10_2 = _zz_PerformanceCounterPlugin_logic_events_sums_10[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_11_2 = _zz_PerformanceCounterPlugin_logic_events_sums_11[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_12_2 = _zz_PerformanceCounterPlugin_logic_events_sums_12[0];
  assign _zz_PerformanceCounterPlugin_logic_events_sums_13_2 = _zz_PerformanceCounterPlugin_logic_events_sums_13[0];
  assign _zz_WhiteboxerPlugin_logic_perf_candidatesCount_1 = DispatchPlugin_logic_candidates_0_ctx_valid;
  assign _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1 = decode_ctrls_1_up_LANE_SEL_0;
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_1 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[9];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_2 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[10];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_3 = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[11],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[12],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[13],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[14],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[15],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[16],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[17],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[18],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[19],{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_4,{_zz_early0_BarrelShifterPlugin_logic_shift_reversed_5,_zz_early0_BarrelShifterPlugin_logic_shift_reversed_6}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_4 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[20];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_5 = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[21];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_reversed_6 = {execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[22],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[23],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[24],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[25],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[26],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[27],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[28],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[29],{execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[30],execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_1 = early0_BarrelShifterPlugin_logic_shift_shifted[9];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_2 = early0_BarrelShifterPlugin_logic_shift_shifted[10];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_3 = {early0_BarrelShifterPlugin_logic_shift_shifted[11],{early0_BarrelShifterPlugin_logic_shift_shifted[12],{early0_BarrelShifterPlugin_logic_shift_shifted[13],{early0_BarrelShifterPlugin_logic_shift_shifted[14],{early0_BarrelShifterPlugin_logic_shift_shifted[15],{early0_BarrelShifterPlugin_logic_shift_shifted[16],{early0_BarrelShifterPlugin_logic_shift_shifted[17],{early0_BarrelShifterPlugin_logic_shift_shifted[18],{early0_BarrelShifterPlugin_logic_shift_shifted[19],{_zz_early0_BarrelShifterPlugin_logic_shift_patched_4,{_zz_early0_BarrelShifterPlugin_logic_shift_patched_5,_zz_early0_BarrelShifterPlugin_logic_shift_patched_6}}}}}}}}}}};
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_4 = early0_BarrelShifterPlugin_logic_shift_shifted[20];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_5 = early0_BarrelShifterPlugin_logic_shift_shifted[21];
  assign _zz_early0_BarrelShifterPlugin_logic_shift_patched_6 = {early0_BarrelShifterPlugin_logic_shift_shifted[22],{early0_BarrelShifterPlugin_logic_shift_shifted[23],{early0_BarrelShifterPlugin_logic_shift_shifted[24],{early0_BarrelShifterPlugin_logic_shift_shifted[25],{early0_BarrelShifterPlugin_logic_shift_shifted[26],{early0_BarrelShifterPlugin_logic_shift_shifted[27],{early0_BarrelShifterPlugin_logic_shift_shifted[28],{early0_BarrelShifterPlugin_logic_shift_shifted[29],{early0_BarrelShifterPlugin_logic_shift_shifted[30],early0_BarrelShifterPlugin_logic_shift_shifted[31]}}}}}}}}};
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1 = _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[6];
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2 = _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[7];
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_3 = {_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[8],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[9],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[10],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[11],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[12],_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[13]}}}}};
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0_1 = 32'h08002054;
  assign _zz_decode_ctrls_1_down_RS2_ENABLE_0_2 = 32'h10002054;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_1 = 32'h00002008;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_2 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000050);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_3 = 32'h00000010;
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000000c) == 32'h00000004);
  assign _zz_decode_ctrls_1_down_RD_ENABLE_0_5 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000028) == 32'h0);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0 = 32'h0000007f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_1 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000107f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_2 = 32'h00001073;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_3 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000207f) == 32'h00002073);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_4 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000407f) == 32'h00004063);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_5 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000207f) == 32'h00002013),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000107f) == 32'h00000013),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_6) == 32'h00000023),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_7 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_8),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_9,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_10,_zz_decode_ctrls_1_down_Decode_LEGAL_0_11}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_6 = 32'h0000603f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_7 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000207f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_8 = 32'h00000003;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_9 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000505f) == 32'h00000003);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_10 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000707b) == 32'h00000063);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_11 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000607f) == 32'h0000000f),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h1800707f) == 32'h0000202f),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_12) == 32'h00000033),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_13 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_14),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_15,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_16,_zz_decode_ctrls_1_down_Decode_LEGAL_0_17}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_12 = 32'hfc00007f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_13 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'he800707f);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_14 = 32'h0800202f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_15 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfc00305f) == 32'h00001013);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_16 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbc00707f) == 32'h00005013);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_17 = {((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbe00707f) == 32'h00005033),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hbe00707f) == 32'h00000033),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0_18) == 32'h1000202f),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_19 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_20),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_21,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_22,_zz_decode_ctrls_1_down_Decode_LEGAL_0_23}}}}}};
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_18 = 32'hf9f0707f;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_19 = (decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hfe007fff);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_20 = 32'h12000073;
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_21 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hdfffffff) == 32'h10200073);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_22 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffefffff) == 32'h00000073);
  assign _zz_decode_ctrls_1_down_Decode_LEGAL_0_23 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'hffffffff) == 32'h10500073);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_1 = 12'ha00;
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_2 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h802) == 12'h002);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_3 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h042) == 12'h0);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_4 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h080) == 12'h080);
  assign _zz_CsrRamPlugin_csrMapper_ramAddress_5 = ((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'h003) == 12'h001);
  assign _zz_GSharePlugin_logic_onLearn_hash_1 = _zz_GSharePlugin_logic_onLearn_hash[6];
  assign _zz_GSharePlugin_logic_onLearn_hash_2 = _zz_GSharePlugin_logic_onLearn_hash[7];
  assign _zz_GSharePlugin_logic_onLearn_hash_3 = {_zz_GSharePlugin_logic_onLearn_hash[8],{_zz_GSharePlugin_logic_onLearn_hash[9],{_zz_GSharePlugin_logic_onLearn_hash[10],{_zz_GSharePlugin_logic_onLearn_hash[11],{_zz_GSharePlugin_logic_onLearn_hash[12],_zz_GSharePlugin_logic_onLearn_hash[13]}}}}};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception}};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception}};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception}};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3 = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception}};
  assign _zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_4 = TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_exception;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated = execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_1 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_2 = execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_3 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_4 = execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_5 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_6 = execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_7 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[21 : 0];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated = fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated_1 = fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0];
  assign _zz_fetch_logic_flushes_0_doIt = 1'b1;
  assign _zz_fetch_logic_flushes_0_doIt_1 = 1'b0;
  assign _zz_fetch_logic_flushes_0_doIt_2 = (1'b1 && BtbPlugin_logic_flushPort_payload_self);
  assign _zz_COMB_CSR_ = 12'hc1f;
  assign _zz_COMB_CSR__1 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1f);
  assign _zz_COMB_CSR__2 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h73e);
  assign _zz_COMB_CSR__3 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc9e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb9e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__4),{_zz_COMB_CSR__5,{_zz_COMB_CSR__6,_zz_COMB_CSR__7}}}}}}}};
  assign _zz_COMB_CSR__4 = 12'h73d;
  assign _zz_COMB_CSR__5 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc9d);
  assign _zz_COMB_CSR__6 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb9d);
  assign _zz_COMB_CSR__7 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33d),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1d),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1d),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h73c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc9c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__8),{_zz_COMB_CSR__9,{_zz_COMB_CSR__10,_zz_COMB_CSR__11}}}}}}}};
  assign _zz_COMB_CSR__8 = 12'hb9c;
  assign _zz_COMB_CSR__9 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33c);
  assign _zz_COMB_CSR__10 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1c);
  assign _zz_COMB_CSR__11 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h73b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc9b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb9b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__12),{_zz_COMB_CSR__13,{_zz_COMB_CSR__14,_zz_COMB_CSR__15}}}}}}}};
  assign _zz_COMB_CSR__12 = 12'hc1b;
  assign _zz_COMB_CSR__13 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1b);
  assign _zz_COMB_CSR__14 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h73a);
  assign _zz_COMB_CSR__15 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc9a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb9a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc1a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb1a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__16),{_zz_COMB_CSR__17,{_zz_COMB_CSR__18,_zz_COMB_CSR__19}}}}}}}};
  assign _zz_COMB_CSR__16 = 12'h739;
  assign _zz_COMB_CSR__17 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc99);
  assign _zz_COMB_CSR__18 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb99);
  assign _zz_COMB_CSR__19 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h339),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc19),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb19),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h738),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc98),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__20),{_zz_COMB_CSR__21,{_zz_COMB_CSR__22,_zz_COMB_CSR__23}}}}}}}};
  assign _zz_COMB_CSR__20 = 12'hb98;
  assign _zz_COMB_CSR__21 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h338);
  assign _zz_COMB_CSR__22 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc18);
  assign _zz_COMB_CSR__23 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb18),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h737),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc97),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb97),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h337),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__24),{_zz_COMB_CSR__25,{_zz_COMB_CSR__26,_zz_COMB_CSR__27}}}}}}}};
  assign _zz_COMB_CSR__24 = 12'hc17;
  assign _zz_COMB_CSR__25 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb17);
  assign _zz_COMB_CSR__26 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h736);
  assign _zz_COMB_CSR__27 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc96),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb96),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h336),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc16),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb16),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__28),{_zz_COMB_CSR__29,{_zz_COMB_CSR__30,_zz_COMB_CSR__31}}}}}}}};
  assign _zz_COMB_CSR__28 = 12'h735;
  assign _zz_COMB_CSR__29 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc95);
  assign _zz_COMB_CSR__30 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb95);
  assign _zz_COMB_CSR__31 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h335),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc15),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb15),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h734),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc94),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__32),{_zz_COMB_CSR__33,{_zz_COMB_CSR__34,_zz_COMB_CSR__35}}}}}}}};
  assign _zz_COMB_CSR__32 = 12'hb94;
  assign _zz_COMB_CSR__33 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h334);
  assign _zz_COMB_CSR__34 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc14);
  assign _zz_COMB_CSR__35 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb14),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h733),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc93),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb93),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h333),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__36),{_zz_COMB_CSR__37,{_zz_COMB_CSR__38,_zz_COMB_CSR__39}}}}}}}};
  assign _zz_COMB_CSR__36 = 12'hc13;
  assign _zz_COMB_CSR__37 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb13);
  assign _zz_COMB_CSR__38 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h732);
  assign _zz_COMB_CSR__39 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc92),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb92),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h332),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc12),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb12),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__40),{_zz_COMB_CSR__41,{_zz_COMB_CSR__42,_zz_COMB_CSR__43}}}}}}}};
  assign _zz_COMB_CSR__40 = 12'h731;
  assign _zz_COMB_CSR__41 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc91);
  assign _zz_COMB_CSR__42 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb91);
  assign _zz_COMB_CSR__43 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h331),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc11),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb11),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h730),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc90),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__44),{_zz_COMB_CSR__45,{_zz_COMB_CSR__46,_zz_COMB_CSR__47}}}}}}}};
  assign _zz_COMB_CSR__44 = 12'hb90;
  assign _zz_COMB_CSR__45 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h330);
  assign _zz_COMB_CSR__46 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc10);
  assign _zz_COMB_CSR__47 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb10),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h72f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc8f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb8f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__48),{_zz_COMB_CSR__49,{_zz_COMB_CSR__50,_zz_COMB_CSR__51}}}}}}}};
  assign _zz_COMB_CSR__48 = 12'hc0f;
  assign _zz_COMB_CSR__49 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0f);
  assign _zz_COMB_CSR__50 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h72e);
  assign _zz_COMB_CSR__51 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc8e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb8e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0e),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__52),{_zz_COMB_CSR__53,{_zz_COMB_CSR__54,_zz_COMB_CSR__55}}}}}}}};
  assign _zz_COMB_CSR__52 = 12'h72d;
  assign _zz_COMB_CSR__53 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc8d);
  assign _zz_COMB_CSR__54 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb8d);
  assign _zz_COMB_CSR__55 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32d),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0d),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0d),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h72c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc8c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__56),{_zz_COMB_CSR__57,{_zz_COMB_CSR__58,_zz_COMB_CSR__59}}}}}}}};
  assign _zz_COMB_CSR__56 = 12'hb8c;
  assign _zz_COMB_CSR__57 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32c);
  assign _zz_COMB_CSR__58 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0c);
  assign _zz_COMB_CSR__59 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0c),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h72b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc8b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb8b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32b),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__60),{_zz_COMB_CSR__61,{_zz_COMB_CSR__62,_zz_COMB_CSR__63}}}}}}}};
  assign _zz_COMB_CSR__60 = 12'hc0b;
  assign _zz_COMB_CSR__61 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0b);
  assign _zz_COMB_CSR__62 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h72a);
  assign _zz_COMB_CSR__63 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc8a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb8a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h32a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc0a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb0a),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__64),{_zz_COMB_CSR__65,{_zz_COMB_CSR__66,_zz_COMB_CSR__67}}}}}}}};
  assign _zz_COMB_CSR__64 = 12'h729;
  assign _zz_COMB_CSR__65 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc89);
  assign _zz_COMB_CSR__66 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb89);
  assign _zz_COMB_CSR__67 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h329),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc09),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb09),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h728),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc88),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__68),{_zz_COMB_CSR__69,{_zz_COMB_CSR__70,_zz_COMB_CSR__71}}}}}}}};
  assign _zz_COMB_CSR__68 = 12'hb88;
  assign _zz_COMB_CSR__69 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h328);
  assign _zz_COMB_CSR__70 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc08);
  assign _zz_COMB_CSR__71 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb08),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h727),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc87),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb87),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h327),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__72),{_zz_COMB_CSR__73,{_zz_COMB_CSR__74,_zz_COMB_CSR__75}}}}}}}};
  assign _zz_COMB_CSR__72 = 12'hc07;
  assign _zz_COMB_CSR__73 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb07);
  assign _zz_COMB_CSR__74 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h726);
  assign _zz_COMB_CSR__75 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc86),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb86),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h326),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc06),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb06),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__76),{_zz_COMB_CSR__77,{_zz_COMB_CSR__78,_zz_COMB_CSR__79}}}}}}}};
  assign _zz_COMB_CSR__76 = 12'h725;
  assign _zz_COMB_CSR__77 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc85);
  assign _zz_COMB_CSR__78 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb85);
  assign _zz_COMB_CSR__79 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h325),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc05),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb05),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h724),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc84),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR__80),{_zz_COMB_CSR__81,{_zz_COMB_CSR__82,_zz_COMB_CSR__83}}}}}}}};
  assign _zz_COMB_CSR__80 = 12'hb84;
  assign _zz_COMB_CSR__81 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h324);
  assign _zz_COMB_CSR__82 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc04);
  assign _zz_COMB_CSR__83 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb04),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h723),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc83),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb83),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h323),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc03),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb03)}}}}}};
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter = 12'hc00;
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_1 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb00);
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_2 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h140);
  assign _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_3 = {(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h141),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h143),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h105),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h340),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h341),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h343),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h305)}}}}}};
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter = 12'hc00;
  assign _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_1 = 12'hb00;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented = COMB_CSR_3073;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_1 = {COMB_CSR_324,{COMB_CSR_260,{COMB_CSR_322,{COMB_CSR_771,{COMB_CSR_770,{COMB_CSR_772,{COMB_CSR_836,{COMB_CSR_834,{COMB_CSR_769,{COMB_CSR_3860,{_zz_CsrAccessPlugin_logic_fsm_inject_implemented_2,_zz_CsrAccessPlugin_logic_fsm_inject_implemented_3}}}}}}}}}}};
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_2 = COMB_CSR_3859;
  assign _zz_CsrAccessPlugin_logic_fsm_inject_implemented_3 = {COMB_CSR_3858,{COMB_CSR_3857,{COMB_CSR_1954,{COMB_CSR_1953,{COMB_CSR_1952,{COMB_CSR_3008,{COMB_CSR_384,{COMB_CSR_256,COMB_CSR_768}}}}}}}};
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_59);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_64 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_65 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_70);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_74 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_75 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_80);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_85 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_86 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_91);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_96 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_97 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_102);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_107 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_108 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_113);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_118 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_119 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_123);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_127 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_128 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_133);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_138 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_139 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_144);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_149 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_150 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_155);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_160 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_161 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_166);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_171 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_172 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_177);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_180 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_181 ? _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_182 : _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_183);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_196 = (CsrRamPlugin_csrMapper_withRead ? CsrRamPlugin_csrMapper_read_data : _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_197);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_21 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_22 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_24);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_26 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_27 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_29);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_32 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_33 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_34);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_36 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_37 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_38);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_41 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_42 | 32'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_44 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_45 | 32'h0);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_48 = (32'h0 | ((when_CsrService_l198 && REG_CSR_769) ? 32'h40141101 : 32'h0));
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_49 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_50 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_52);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_55 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_56 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_58);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_59 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_60 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_62);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_65 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_66 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_68);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_70 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_71 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_73);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_75 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_76 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_78);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_80 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_81 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_83);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_86 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_87 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_89);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_91 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_92 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_94);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_97 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_98 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_100);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_102 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_103 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_105);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_108 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_109 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_111);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_113 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_114 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_116);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_119 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_120 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_122);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_123 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_124 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_126);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_128 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_129 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_131);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_133 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_134 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_136);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_139 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_140 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_142);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_144 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_145 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_147);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_150 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_151 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_153);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_155 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_156 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_158);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_161 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_162 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_164);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_166 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_167 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_169);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_172 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_173 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_175);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_177 = (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_178 | ((when_CsrService_l198 && REG_CSR_3073) ? PrivilegedPlugin_logic_rdtime[31 : 0] : 32'h0));
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_181 = (when_CsrService_l198 && REG_CSR_3201);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_182 = PrivilegedPlugin_logic_rdtime[63 : 32];
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_183 = 32'h0;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_197 = 32'h0;
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault = 32'hfffff000;
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault_1 = 32'hfffff800;
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_fault = 32'hffff0000;
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_fault_1 = (LsuPlugin_pmaBuilder_l1_addressBits & 32'hfffff000);
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_fault_2 = 32'h10000000;
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_fault_3 = (LsuPlugin_pmaBuilder_l1_addressBits & 32'hfffff800);
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_fault_4 = 32'h10001000;
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault = 32'hffc00000;
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_1 = (LsuPlugin_pmaBuilder_io_addressBits & 32'hfffe0000);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_2 = 32'hf0000000;
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_3 = ((LsuPlugin_pmaBuilder_io_addressBits & 32'hffff0000) == 32'h0);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_4 = ((LsuPlugin_pmaBuilder_io_addressBits & 32'hfffff000) == 32'h10000000);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_fault_5 = ((LsuPlugin_pmaBuilder_io_addressBits & 32'hfffff800) == 32'h10001000);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_3 = (execute_lane0_logic_decoding_decodingBits & 32'h00000050);
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_4 = 32'h00000010;
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_5 = _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0;
  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_6 = _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0;
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = 32'h00002020;
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_1 = (execute_lane0_logic_decoding_decodingBits & 32'h08002000);
  assign _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_2 = 32'h00002000;
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2 = 32'h02001000;
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_1 = 32'h10201000;
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_2 = (execute_lane0_logic_decoding_decodingBits & 32'h12400000);
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_3 = 32'h10000000;
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_4 = ((execute_lane0_logic_decoding_decodingBits & 32'h10100000) == 32'h00100000);
  assign _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_5 = ((execute_lane0_logic_decoding_decodingBits & 32'h12200000) == 32'h10000000);
  assign _zz_when_ExecuteLanePlugin_l306_2 = 1'b1;
  always @(posedge litex_clk) begin
    if(_zz_10) begin
      FetchL1Plugin_logic_banks_0_mem[FetchL1Plugin_logic_banks_0_write_payload_address] <= FetchL1Plugin_logic_banks_0_write_payload_data;
    end
  end

  always @(posedge litex_clk) begin
    if(FetchL1Plugin_logic_banks_0_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_0_mem_spinal_port1 <= FetchL1Plugin_logic_banks_0_mem[FetchL1Plugin_logic_banks_0_read_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_9) begin
      FetchL1Plugin_logic_banks_1_mem[FetchL1Plugin_logic_banks_1_write_payload_address] <= FetchL1Plugin_logic_banks_1_write_payload_data;
    end
  end

  always @(posedge litex_clk) begin
    if(FetchL1Plugin_logic_banks_1_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_1_mem_spinal_port1 <= FetchL1Plugin_logic_banks_1_mem[FetchL1Plugin_logic_banks_1_read_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_8) begin
      FetchL1Plugin_logic_banks_2_mem[FetchL1Plugin_logic_banks_2_write_payload_address] <= FetchL1Plugin_logic_banks_2_write_payload_data;
    end
  end

  always @(posedge litex_clk) begin
    if(FetchL1Plugin_logic_banks_2_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_2_mem_spinal_port1 <= FetchL1Plugin_logic_banks_2_mem[FetchL1Plugin_logic_banks_2_read_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_7) begin
      FetchL1Plugin_logic_banks_3_mem[FetchL1Plugin_logic_banks_3_write_payload_address] <= FetchL1Plugin_logic_banks_3_write_payload_data;
    end
  end

  always @(posedge litex_clk) begin
    if(FetchL1Plugin_logic_banks_3_read_cmd_valid) begin
      FetchL1Plugin_logic_banks_3_mem_spinal_port1 <= FetchL1Plugin_logic_banks_3_mem[FetchL1Plugin_logic_banks_3_read_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_FetchL1Plugin_logic_ways_0_mem_port_1) begin
      FetchL1Plugin_logic_ways_0_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_0_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(FetchL1Plugin_logic_ways_0_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_0_mem_spinal_port1 <= FetchL1Plugin_logic_ways_0_mem[FetchL1Plugin_logic_ways_0_read_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_FetchL1Plugin_logic_ways_1_mem_port_1) begin
      FetchL1Plugin_logic_ways_1_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_1_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(FetchL1Plugin_logic_ways_1_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_1_mem_spinal_port1 <= FetchL1Plugin_logic_ways_1_mem[FetchL1Plugin_logic_ways_1_read_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_FetchL1Plugin_logic_ways_2_mem_port_1) begin
      FetchL1Plugin_logic_ways_2_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_2_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(FetchL1Plugin_logic_ways_2_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_2_mem_spinal_port1 <= FetchL1Plugin_logic_ways_2_mem[FetchL1Plugin_logic_ways_2_read_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_FetchL1Plugin_logic_ways_3_mem_port_1) begin
      FetchL1Plugin_logic_ways_3_mem[FetchL1Plugin_logic_waysWrite_address] <= _zz_FetchL1Plugin_logic_ways_3_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(FetchL1Plugin_logic_ways_3_read_cmd_valid) begin
      FetchL1Plugin_logic_ways_3_mem_spinal_port1 <= FetchL1Plugin_logic_ways_3_mem[FetchL1Plugin_logic_ways_3_read_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_6) begin
      FetchL1Plugin_logic_plru_mem[FetchL1Plugin_logic_plru_write_payload_address] <= _zz_FetchL1Plugin_logic_plru_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(FetchL1Plugin_logic_plru_read_cmd_valid) begin
      FetchL1Plugin_logic_plru_mem_spinal_port1 <= FetchL1Plugin_logic_plru_mem[FetchL1Plugin_logic_plru_read_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_5) begin
      GSharePlugin_logic_mem_counter[GSharePlugin_logic_mem_write_payload_address] <= _zz_GSharePlugin_logic_mem_counter_port;
    end
  end

  always @(posedge litex_clk) begin
    if(fetch_logic_ctrls_0_down_isReady) begin
      GSharePlugin_logic_mem_counter_spinal_port1 <= GSharePlugin_logic_mem_counter[fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH];
    end
  end

  always @(posedge litex_clk) begin
    if(BtbPlugin_logic_memDp_wp_payload_mask[0] && BtbPlugin_logic_memDp_wp_valid) begin
      BtbPlugin_logic_mem[BtbPlugin_logic_memDp_wp_payload_address] <= _zz_BtbPlugin_logic_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(BtbPlugin_logic_memDp_rp_cmd_valid) begin
      BtbPlugin_logic_mem_spinal_port1 <= BtbPlugin_logic_mem[BtbPlugin_logic_memDp_rp_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_LsuL1Plugin_logic_ways_0_mem_port_1) begin
      LsuL1Plugin_logic_ways_0_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_0_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_0_mem_spinal_port1 <= LsuL1Plugin_logic_ways_0_mem[LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_LsuL1Plugin_logic_ways_1_mem_port_1) begin
      LsuL1Plugin_logic_ways_1_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_1_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_1_mem_spinal_port1 <= LsuL1Plugin_logic_ways_1_mem[LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_LsuL1Plugin_logic_ways_2_mem_port_1) begin
      LsuL1Plugin_logic_ways_2_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_2_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(LsuL1Plugin_logic_ways_2_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_2_mem_spinal_port1 <= LsuL1Plugin_logic_ways_2_mem[LsuL1Plugin_logic_ways_2_lsuRead_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_LsuL1Plugin_logic_ways_3_mem_port_1) begin
      LsuL1Plugin_logic_ways_3_mem[LsuL1Plugin_logic_waysWrite_address] <= _zz_LsuL1Plugin_logic_ways_3_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(LsuL1Plugin_logic_ways_3_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_ways_3_mem_spinal_port1 <= LsuL1Plugin_logic_ways_3_mem[LsuL1Plugin_logic_ways_3_lsuRead_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_4) begin
      LsuL1Plugin_logic_shared_mem[LsuL1Plugin_logic_shared_write_payload_address] <= _zz_LsuL1Plugin_logic_shared_mem_port;
    end
  end

  always @(posedge litex_clk) begin
    if(LsuL1Plugin_logic_shared_lsuRead_cmd_valid) begin
      LsuL1Plugin_logic_shared_mem_spinal_port1 <= LsuL1Plugin_logic_shared_mem[LsuL1Plugin_logic_shared_lsuRead_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_3) begin
      LsuL1Plugin_logic_writeback_victimBuffer[_zz_LsuL1Plugin_logic_writeback_victimBuffer_port] <= LsuL1Plugin_logic_writeback_read_readedData;
    end
  end

  always @(posedge litex_clk) begin
    if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
      LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1 <= LsuL1Plugin_logic_writeback_victimBuffer[_zz_LsuL1Plugin_logic_writeback_write_word];
    end
  end

  always @(posedge litex_clk) begin
    if(_zz_2) begin
      CsrRamPlugin_logic_mem[CsrRamPlugin_logic_writeLogic_port_payload_address] <= CsrRamPlugin_logic_writeLogic_port_payload_data;
    end
  end

  always @(posedge litex_clk) begin
    if(CsrRamPlugin_logic_readLogic_port_cmd_valid) begin
      CsrRamPlugin_logic_mem_spinal_port1 <= CsrRamPlugin_logic_mem[CsrRamPlugin_logic_readLogic_port_cmd_payload];
    end
  end

  DivRadix early0_DivPlugin_logic_processing_div (
    .io_flush                  (execute_ctrl2_down_isReady                                       ), //i
    .io_cmd_valid              (early0_DivPlugin_logic_processing_div_io_cmd_valid               ), //i
    .io_cmd_ready              (early0_DivPlugin_logic_processing_div_io_cmd_ready               ), //o
    .io_cmd_payload_a          (early0_DivPlugin_logic_processing_a[31:0]                        ), //i
    .io_cmd_payload_b          (early0_DivPlugin_logic_processing_b[31:0]                        ), //i
    .io_cmd_payload_normalized (1'b0                                                             ), //i
    .io_cmd_payload_iterations (5'bxxxxx                                                         ), //i
    .io_rsp_valid              (early0_DivPlugin_logic_processing_div_io_rsp_valid               ), //o
    .io_rsp_ready              (1'b0                                                             ), //i
    .io_rsp_payload_result     (early0_DivPlugin_logic_processing_div_io_rsp_payload_result[31:0]), //o
    .io_rsp_payload_remain     (early0_DivPlugin_logic_processing_div_io_rsp_payload_remain[31:0]), //o
    .litex_clk                 (litex_clk                                                        ), //i
    .cpuResetCtrl_reset        (cpuResetCtrl_reset                                               )  //i
  );
  StreamFifoLowLatency CfuPlugin_logic_onJoin_busRspStream_fifo (
    .io_push_valid             (CfuPlugin_logic_onJoin_busRspStream_valid                              ), //i
    .io_push_ready             (CfuPlugin_logic_onJoin_busRspStream_fifo_io_push_ready                 ), //o
    .io_push_payload_outputs_0 (CfuPlugin_logic_onJoin_busRspStream_payload_outputs_0[31:0]            ), //i
    .io_pop_valid              (CfuPlugin_logic_onJoin_busRspStream_fifo_io_pop_valid                  ), //o
    .io_pop_ready              (CfuPlugin_logic_onJoin_busRspStream_fifo_io_pop_ready                  ), //i
    .io_pop_payload_outputs_0  (CfuPlugin_logic_onJoin_busRspStream_fifo_io_pop_payload_outputs_0[31:0]), //o
    .io_flush                  (1'b0                                                                   ), //i
    .io_occupancy              (CfuPlugin_logic_onJoin_busRspStream_fifo_io_occupancy[1:0]             ), //o
    .io_availability           (CfuPlugin_logic_onJoin_busRspStream_fifo_io_availability[1:0]          ), //o
    .litex_clk                 (litex_clk                                                              ), //i
    .cpuResetCtrl_reset        (cpuResetCtrl_reset                                                     )  //i
  );
  StreamArbiter LsuPlugin_logic_flusher_arbiter (
    .io_inputs_0_valid  (TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid     ), //i
    .io_inputs_0_ready  (LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready), //o
    .io_output_valid    (LsuPlugin_logic_flusher_arbiter_io_output_valid  ), //o
    .io_output_ready    (LsuPlugin_logic_flusher_arbiter_io_output_ready  ), //i
    .io_chosenOH        (LsuPlugin_logic_flusher_arbiter_io_chosenOH      ), //o
    .litex_clk          (litex_clk                                        ), //i
    .cpuResetCtrl_reset (cpuResetCtrl_reset                               )  //i
  );
  StreamArbiter_1 streamArbiter_10 (
    .io_inputs_0_valid                                     (LearnPlugin_logic_buffered_0_valid                                         ), //i
    .io_inputs_0_ready                                     (streamArbiter_10_io_inputs_0_ready                                         ), //o
    .io_inputs_0_payload_pcOnLastSlice                     (LearnPlugin_logic_buffered_0_payload_pcOnLastSlice[31:0]                   ), //i
    .io_inputs_0_payload_pcTarget                          (LearnPlugin_logic_buffered_0_payload_pcTarget[31:0]                        ), //i
    .io_inputs_0_payload_taken                             (LearnPlugin_logic_buffered_0_payload_taken                                 ), //i
    .io_inputs_0_payload_isBranch                          (LearnPlugin_logic_buffered_0_payload_isBranch                              ), //i
    .io_inputs_0_payload_isPush                            (LearnPlugin_logic_buffered_0_payload_isPush                                ), //i
    .io_inputs_0_payload_isPop                             (LearnPlugin_logic_buffered_0_payload_isPop                                 ), //i
    .io_inputs_0_payload_wasWrong                          (LearnPlugin_logic_buffered_0_payload_wasWrong                              ), //i
    .io_inputs_0_payload_badPredictedTarget                (LearnPlugin_logic_buffered_0_payload_badPredictedTarget                    ), //i
    .io_inputs_0_payload_history                           (LearnPlugin_logic_buffered_0_payload_history[11:0]                         ), //i
    .io_inputs_0_payload_uopId                             (LearnPlugin_logic_buffered_0_payload_uopId[15:0]                           ), //i
    .io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 (LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]), //i
    .io_output_valid                                       (streamArbiter_10_io_output_valid                                           ), //o
    .io_output_ready                                       (LearnPlugin_logic_arbitrated_ready                                         ), //i
    .io_output_payload_pcOnLastSlice                       (streamArbiter_10_io_output_payload_pcOnLastSlice[31:0]                     ), //o
    .io_output_payload_pcTarget                            (streamArbiter_10_io_output_payload_pcTarget[31:0]                          ), //o
    .io_output_payload_taken                               (streamArbiter_10_io_output_payload_taken                                   ), //o
    .io_output_payload_isBranch                            (streamArbiter_10_io_output_payload_isBranch                                ), //o
    .io_output_payload_isPush                              (streamArbiter_10_io_output_payload_isPush                                  ), //o
    .io_output_payload_isPop                               (streamArbiter_10_io_output_payload_isPop                                   ), //o
    .io_output_payload_wasWrong                            (streamArbiter_10_io_output_payload_wasWrong                                ), //o
    .io_output_payload_badPredictedTarget                  (streamArbiter_10_io_output_payload_badPredictedTarget                      ), //o
    .io_output_payload_history                             (streamArbiter_10_io_output_payload_history[11:0]                           ), //o
    .io_output_payload_uopId                               (streamArbiter_10_io_output_payload_uopId[15:0]                             ), //o
    .io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0   (streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1:0]  ), //o
    .io_chosenOH                                           (streamArbiter_10_io_chosenOH                                               ), //o
    .litex_clk                                             (litex_clk                                                                  ), //i
    .cpuResetCtrl_reset                                    (cpuResetCtrl_reset                                                         )  //i
  );
  StreamArbiter_2 LsuPlugin_logic_onAddress0_arbiter (
    .io_inputs_0_valid              (LsuPlugin_logic_onAddress0_ls_port_valid                          ), //i
    .io_inputs_0_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready              ), //o
    .io_inputs_0_payload_op         (LsuPlugin_logic_onAddress0_ls_port_payload_op[2:0]                ), //i
    .io_inputs_0_payload_address    (LsuPlugin_logic_onAddress0_ls_port_payload_address[31:0]          ), //i
    .io_inputs_0_payload_size       (LsuPlugin_logic_onAddress0_ls_port_payload_size[1:0]              ), //i
    .io_inputs_0_payload_load       (LsuPlugin_logic_onAddress0_ls_port_payload_load                   ), //i
    .io_inputs_0_payload_store      (LsuPlugin_logic_onAddress0_ls_port_payload_store                  ), //i
    .io_inputs_0_payload_atomic     (LsuPlugin_logic_onAddress0_ls_port_payload_atomic                 ), //i
    .io_inputs_0_payload_clean      (LsuPlugin_logic_onAddress0_ls_port_payload_clean                  ), //i
    .io_inputs_0_payload_invalidate (LsuPlugin_logic_onAddress0_ls_port_payload_invalidate             ), //i
    .io_inputs_0_payload_storeId    (LsuPlugin_logic_onAddress0_ls_port_payload_storeId[11:0]          ), //i
    .io_inputs_1_valid              (LsuPlugin_logic_onAddress0_access_port_valid                      ), //i
    .io_inputs_1_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready              ), //o
    .io_inputs_1_payload_op         (LsuPlugin_logic_onAddress0_access_port_payload_op[2:0]            ), //i
    .io_inputs_1_payload_address    (LsuPlugin_logic_onAddress0_access_port_payload_address[31:0]      ), //i
    .io_inputs_1_payload_size       (LsuPlugin_logic_onAddress0_access_port_payload_size[1:0]          ), //i
    .io_inputs_1_payload_load       (LsuPlugin_logic_onAddress0_access_port_payload_load               ), //i
    .io_inputs_1_payload_store      (LsuPlugin_logic_onAddress0_access_port_payload_store              ), //i
    .io_inputs_1_payload_atomic     (LsuPlugin_logic_onAddress0_access_port_payload_atomic             ), //i
    .io_inputs_1_payload_clean      (LsuPlugin_logic_onAddress0_access_port_payload_clean              ), //i
    .io_inputs_1_payload_invalidate (LsuPlugin_logic_onAddress0_access_port_payload_invalidate         ), //i
    .io_inputs_1_payload_storeId    (LsuPlugin_logic_onAddress0_access_port_payload_storeId[11:0]      ), //i
    .io_inputs_2_valid              (LsuPlugin_logic_onAddress0_flush_port_valid                       ), //i
    .io_inputs_2_ready              (LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready              ), //o
    .io_inputs_2_payload_op         (LsuPlugin_logic_onAddress0_flush_port_payload_op[2:0]             ), //i
    .io_inputs_2_payload_address    (LsuPlugin_logic_onAddress0_flush_port_payload_address[31:0]       ), //i
    .io_inputs_2_payload_size       (LsuPlugin_logic_onAddress0_flush_port_payload_size[1:0]           ), //i
    .io_inputs_2_payload_load       (LsuPlugin_logic_onAddress0_flush_port_payload_load                ), //i
    .io_inputs_2_payload_store      (LsuPlugin_logic_onAddress0_flush_port_payload_store               ), //i
    .io_inputs_2_payload_atomic     (LsuPlugin_logic_onAddress0_flush_port_payload_atomic              ), //i
    .io_inputs_2_payload_clean      (LsuPlugin_logic_onAddress0_flush_port_payload_clean               ), //i
    .io_inputs_2_payload_invalidate (LsuPlugin_logic_onAddress0_flush_port_payload_invalidate          ), //i
    .io_inputs_2_payload_storeId    (LsuPlugin_logic_onAddress0_flush_port_payload_storeId[11:0]       ), //i
    .io_output_valid                (LsuPlugin_logic_onAddress0_arbiter_io_output_valid                ), //o
    .io_output_ready                (LsuPlugin_logic_onAddress0_arbiter_io_output_ready                ), //i
    .io_output_payload_op           (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op[2:0]      ), //o
    .io_output_payload_address      (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address[31:0]), //o
    .io_output_payload_size         (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size[1:0]    ), //o
    .io_output_payload_load         (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load         ), //o
    .io_output_payload_store        (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store        ), //o
    .io_output_payload_atomic       (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic       ), //o
    .io_output_payload_clean        (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_clean        ), //o
    .io_output_payload_invalidate   (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_invalidate   ), //o
    .io_output_payload_storeId      (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId[11:0]), //o
    .io_chosen                      (LsuPlugin_logic_onAddress0_arbiter_io_chosen[1:0]                 ), //o
    .io_chosenOH                    (LsuPlugin_logic_onAddress0_arbiter_io_chosenOH[2:0]               ), //o
    .litex_clk                      (litex_clk                                                         ), //i
    .cpuResetCtrl_reset             (cpuResetCtrl_reset                                                )  //i
  );
  StreamArbiter_3 MmuPlugin_logic_refill_arbiter (
    .io_inputs_0_valid             (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid                ), //i
    .io_inputs_0_ready             (MmuPlugin_logic_refill_arbiter_io_inputs_0_ready                           ), //o
    .io_inputs_0_payload_address   (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_address[31:0]), //i
    .io_inputs_0_payload_storageId (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_storageId    ), //i
    .io_output_valid               (MmuPlugin_logic_refill_arbiter_io_output_valid                             ), //o
    .io_output_ready               (MmuPlugin_logic_refill_arbiter_io_output_ready                             ), //i
    .io_output_payload_address     (MmuPlugin_logic_refill_arbiter_io_output_payload_address[31:0]             ), //o
    .io_output_payload_storageId   (MmuPlugin_logic_refill_arbiter_io_output_payload_storageId                 ), //o
    .io_chosenOH                   (MmuPlugin_logic_refill_arbiter_io_chosenOH                                 ), //o
    .litex_clk                     (litex_clk                                                                  ), //i
    .cpuResetCtrl_reset            (cpuResetCtrl_reset                                                         )  //i
  );
  StreamArbiter_4 MmuPlugin_logic_invalidate_arbiter (
    .io_inputs_0_valid  (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid), //i
    .io_inputs_0_ready  (MmuPlugin_logic_invalidate_arbiter_io_inputs_0_ready           ), //o
    .io_output_valid    (MmuPlugin_logic_invalidate_arbiter_io_output_valid             ), //o
    .io_output_ready    (MmuPlugin_logic_invalidate_arbiter_io_output_ready             ), //i
    .io_chosenOH        (MmuPlugin_logic_invalidate_arbiter_io_chosenOH                 ), //o
    .litex_clk          (litex_clk                                                      ), //i
    .cpuResetCtrl_reset (cpuResetCtrl_reset                                             )  //i
  );
  RegFileMem integer_RegFilePlugin_logic_regfile_fpga (
    .io_writes_0_valid   (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid       ), //i
    .io_writes_0_address (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address[4:0]), //i
    .io_writes_0_data    (integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data[31:0]  ), //i
    .io_writes_0_uopId   (integer_RegFilePlugin_logic_writeMerges_0_bus_uopId[15:0]        ), //i
    .io_reads_0_valid    (execute_lane0_bypasser_integer_RS1_port_valid                    ), //i
    .io_reads_0_address  (execute_lane0_bypasser_integer_RS1_port_address[4:0]             ), //i
    .io_reads_0_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data[31:0]   ), //o
    .io_reads_1_valid    (execute_lane0_bypasser_integer_RS2_port_valid                    ), //i
    .io_reads_1_address  (execute_lane0_bypasser_integer_RS2_port_address[4:0]             ), //i
    .io_reads_1_data     (integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data[31:0]   ), //o
    .litex_clk           (litex_clk                                                        ), //i
    .cpuResetCtrl_reset  (cpuResetCtrl_reset                                               )  //i
  );
  Ram_1w_1ra #(
    .wordCount      (4         ),
    .wordWidth      (30        ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (2         ),
    .wrDataWidth    (30        ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (2         ),
    .rdDataWidth    (30        )
  ) BtbPlugin_logic_ras_mem_stack (
    .clk     (litex_clk                                     ), //i
    .wr_en   (BtbPlugin_logic_ras_mem_stack_wr_en           ), //i
    .wr_mask (1'b1                                          ), //i
    .wr_addr (BtbPlugin_logic_ras_write_payload_address[1:0]), //i
    .wr_data (BtbPlugin_logic_ras_mem_stack_wr_data[29:0]   ), //i
    .rd_addr (BtbPlugin_logic_ras_ptr_pop_aheadValue[1:0]   ), //i
    .rd_data (BtbPlugin_logic_ras_mem_stack_rd_data[29:0]   )  //o
  );
  Ram_1w_1rs #(
    .wordCount      (512       ),
    .wordWidth      (64        ),
    .clockCrossing  (1'b0      ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (9         ),
    .wrDataWidth    (64        ),
    .wrMaskWidth    (8         ),
    .wrMaskEnable   (1'b1      ),
    .rdAddressWidth (9         ),
    .rdDataWidth    (64        ),
    .rdLatency      (1         )
  ) LsuL1Plugin_logic_banks_0_mem (
    .wr_clk    (litex_clk                                           ), //i
    .wr_en     (LsuL1Plugin_logic_banks_0_mem_wr_en                 ), //i
    .wr_mask   (LsuL1Plugin_logic_banks_0_write_payload_mask[7:0]   ), //i
    .wr_addr   (LsuL1Plugin_logic_banks_0_write_payload_address[8:0]), //i
    .wr_data   (LsuL1Plugin_logic_banks_0_write_payload_data[63:0]  ), //i
    .rd_clk    (litex_clk                                           ), //i
    .rd_en     (LsuL1Plugin_logic_banks_0_mem_rd_en                 ), //i
    .rd_addr   (LsuL1Plugin_logic_banks_0_read_cmd_payload[8:0]     ), //i
    .rd_dataEn (1'b1                                                ), //i
    .rd_data   (LsuL1Plugin_logic_banks_0_mem_rd_data[63:0]         )  //o
  );
  Ram_1w_1rs #(
    .wordCount      (512       ),
    .wordWidth      (64        ),
    .clockCrossing  (1'b0      ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (9         ),
    .wrDataWidth    (64        ),
    .wrMaskWidth    (8         ),
    .wrMaskEnable   (1'b1      ),
    .rdAddressWidth (9         ),
    .rdDataWidth    (64        ),
    .rdLatency      (1         )
  ) LsuL1Plugin_logic_banks_1_mem (
    .wr_clk    (litex_clk                                           ), //i
    .wr_en     (LsuL1Plugin_logic_banks_1_mem_wr_en                 ), //i
    .wr_mask   (LsuL1Plugin_logic_banks_1_write_payload_mask[7:0]   ), //i
    .wr_addr   (LsuL1Plugin_logic_banks_1_write_payload_address[8:0]), //i
    .wr_data   (LsuL1Plugin_logic_banks_1_write_payload_data[63:0]  ), //i
    .rd_clk    (litex_clk                                           ), //i
    .rd_en     (LsuL1Plugin_logic_banks_1_mem_rd_en                 ), //i
    .rd_addr   (LsuL1Plugin_logic_banks_1_read_cmd_payload[8:0]     ), //i
    .rd_dataEn (1'b1                                                ), //i
    .rd_data   (LsuL1Plugin_logic_banks_1_mem_rd_data[63:0]         )  //o
  );
  Ram_1w_1rs #(
    .wordCount      (512       ),
    .wordWidth      (64        ),
    .clockCrossing  (1'b0      ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (9         ),
    .wrDataWidth    (64        ),
    .wrMaskWidth    (8         ),
    .wrMaskEnable   (1'b1      ),
    .rdAddressWidth (9         ),
    .rdDataWidth    (64        ),
    .rdLatency      (1         )
  ) LsuL1Plugin_logic_banks_2_mem (
    .wr_clk    (litex_clk                                           ), //i
    .wr_en     (LsuL1Plugin_logic_banks_2_mem_wr_en                 ), //i
    .wr_mask   (LsuL1Plugin_logic_banks_2_write_payload_mask[7:0]   ), //i
    .wr_addr   (LsuL1Plugin_logic_banks_2_write_payload_address[8:0]), //i
    .wr_data   (LsuL1Plugin_logic_banks_2_write_payload_data[63:0]  ), //i
    .rd_clk    (litex_clk                                           ), //i
    .rd_en     (LsuL1Plugin_logic_banks_2_mem_rd_en                 ), //i
    .rd_addr   (LsuL1Plugin_logic_banks_2_read_cmd_payload[8:0]     ), //i
    .rd_dataEn (1'b1                                                ), //i
    .rd_data   (LsuL1Plugin_logic_banks_2_mem_rd_data[63:0]         )  //o
  );
  Ram_1w_1rs #(
    .wordCount      (512       ),
    .wordWidth      (64        ),
    .clockCrossing  (1'b0      ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (9         ),
    .wrDataWidth    (64        ),
    .wrMaskWidth    (8         ),
    .wrMaskEnable   (1'b1      ),
    .rdAddressWidth (9         ),
    .rdDataWidth    (64        ),
    .rdLatency      (1         )
  ) LsuL1Plugin_logic_banks_3_mem (
    .wr_clk    (litex_clk                                           ), //i
    .wr_en     (LsuL1Plugin_logic_banks_3_mem_wr_en                 ), //i
    .wr_mask   (LsuL1Plugin_logic_banks_3_write_payload_mask[7:0]   ), //i
    .wr_addr   (LsuL1Plugin_logic_banks_3_write_payload_address[8:0]), //i
    .wr_data   (LsuL1Plugin_logic_banks_3_write_payload_data[63:0]  ), //i
    .rd_clk    (litex_clk                                           ), //i
    .rd_en     (LsuL1Plugin_logic_banks_3_mem_rd_en                 ), //i
    .rd_addr   (LsuL1Plugin_logic_banks_3_read_cmd_payload[8:0]     ), //i
    .rd_dataEn (1'b1                                                ), //i
    .rd_data   (LsuL1Plugin_logic_banks_3_mem_rd_data[63:0]         )  //o
  );
  Ram_1w_1ra #(
    .wordCount      (32        ),
    .wordWidth      (40        ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (5         ),
    .wrDataWidth    (40        ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (5         ),
    .rdDataWidth    (40        )
  ) FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0 (
    .clk     (litex_clk                                                             ), //i
    .wr_en   (FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_wr_en        ), //i
    .wr_mask (1'b1                                                                  ), //i
    .wr_addr (FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address[4:0]  ), //i
    .wr_data (FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_wr_data[39:0]), //i
    .rd_addr (FetchL1Plugin_logic_translationPort_logic_read_0_readAddress[4:0]     ), //i
    .rd_data (FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_rd_data[39:0])  //o
  );
  Ram_1w_1ra #(
    .wordCount      (32        ),
    .wordWidth      (40        ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (5         ),
    .wrDataWidth    (40        ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (5         ),
    .rdDataWidth    (40        )
  ) FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1 (
    .clk     (litex_clk                                                             ), //i
    .wr_en   (FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_wr_en        ), //i
    .wr_mask (1'b1                                                                  ), //i
    .wr_addr (FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address[4:0]  ), //i
    .wr_data (FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_wr_data[39:0]), //i
    .rd_addr (FetchL1Plugin_logic_translationPort_logic_read_0_readAddress[4:0]     ), //i
    .rd_data (FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_rd_data[39:0])  //o
  );
  Ram_1w_1ra #(
    .wordCount      (32        ),
    .wordWidth      (20        ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (5         ),
    .wrDataWidth    (20        ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (5         ),
    .rdDataWidth    (20        )
  ) FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0 (
    .clk     (litex_clk                                                             ), //i
    .wr_en   (FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_wr_en        ), //i
    .wr_mask (1'b1                                                                  ), //i
    .wr_addr (FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address[4:0]  ), //i
    .wr_data (FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_wr_data[19:0]), //i
    .rd_addr (FetchL1Plugin_logic_translationPort_logic_read_1_readAddress[4:0]     ), //i
    .rd_data (FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_rd_data[19:0])  //o
  );
  Ram_1w_1ra #(
    .wordCount      (32        ),
    .wordWidth      (40        ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (5         ),
    .wrDataWidth    (40        ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (5         ),
    .rdDataWidth    (40        )
  ) LsuPlugin_logic_translationStorage_logic_sl_0_ways_0 (
    .clk     (litex_clk                                                               ), //i
    .wr_en   (LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_wr_en              ), //i
    .wr_mask (1'b1                                                                    ), //i
    .wr_addr (LsuPlugin_logic_translationStorage_logic_sl_0_write_address[4:0]        ), //i
    .wr_data (LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_wr_data[39:0]      ), //i
    .rd_addr (LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress[4:0]), //i
    .rd_data (LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_rd_data[39:0]      )  //o
  );
  Ram_1w_1ra #(
    .wordCount      (32        ),
    .wordWidth      (40        ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (5         ),
    .wrDataWidth    (40        ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (5         ),
    .rdDataWidth    (40        )
  ) LsuPlugin_logic_translationStorage_logic_sl_0_ways_1 (
    .clk     (litex_clk                                                               ), //i
    .wr_en   (LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_wr_en              ), //i
    .wr_mask (1'b1                                                                    ), //i
    .wr_addr (LsuPlugin_logic_translationStorage_logic_sl_0_write_address[4:0]        ), //i
    .wr_data (LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_wr_data[39:0]      ), //i
    .rd_addr (LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress[4:0]), //i
    .rd_data (LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_rd_data[39:0]      )  //o
  );
  Ram_1w_1ra #(
    .wordCount      (32        ),
    .wordWidth      (40        ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (5         ),
    .wrDataWidth    (40        ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (5         ),
    .rdDataWidth    (40        )
  ) LsuPlugin_logic_translationStorage_logic_sl_0_ways_2 (
    .clk     (litex_clk                                                               ), //i
    .wr_en   (LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_wr_en              ), //i
    .wr_mask (1'b1                                                                    ), //i
    .wr_addr (LsuPlugin_logic_translationStorage_logic_sl_0_write_address[4:0]        ), //i
    .wr_data (LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_wr_data[39:0]      ), //i
    .rd_addr (LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress[4:0]), //i
    .rd_data (LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_rd_data[39:0]      )  //o
  );
  Ram_1w_1ra #(
    .wordCount      (32        ),
    .wordWidth      (20        ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (5         ),
    .wrDataWidth    (20        ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (5         ),
    .rdDataWidth    (20        )
  ) LsuPlugin_logic_translationStorage_logic_sl_1_ways_0 (
    .clk     (litex_clk                                                               ), //i
    .wr_en   (LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_wr_en              ), //i
    .wr_mask (1'b1                                                                    ), //i
    .wr_addr (LsuPlugin_logic_translationStorage_logic_sl_1_write_address[4:0]        ), //i
    .wr_data (LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_wr_data[19:0]      ), //i
    .rd_addr (LsuPlugin_logic_onAddress0_translationPort_logic_read_1_readAddress[4:0]), //i
    .rd_data (LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_rd_data[19:0]      )  //o
  );
  always @(*) begin
    case(_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0_1)
      1'b0 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0[31 : 0];
      default : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1_1)
      1'b0 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1[31 : 0];
      default : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2_1)
      1'b0 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_2[31 : 0];
      default : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_2[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3_1)
      1'b0 : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_3[31 : 0];
      default : _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_3[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_commitCount_1)
      1'b0 : _zz_PerformanceCounterPlugin_logic_commitCount = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_commitCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(execute_ctrl2_down_CfuPlugin_logic_CFU_ENCODING_lane0)
      1'b0 : _zz_CfuPlugin_logic_bus_cmd_payload_function_id = CfuPlugin_logic_onFork_functionsIds_0;
      default : _zz_CfuPlugin_logic_bus_cmd_payload_function_id = CfuPlugin_logic_onFork_functionsIds_1;
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way)
      2'b00 : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_0_read_rsp;
      2'b01 : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_1_read_rsp;
      2'b10 : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_2_read_rsp;
      default : _zz_LsuL1Plugin_logic_writeback_read_readedData = LsuL1Plugin_logic_banks_3_read_rsp;
    endcase
  end

  always @(*) begin
    case(_zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0_1)
      1'b0 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0[31 : 0];
      default : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1_1)
      1'b0 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1[31 : 0];
      default : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2_1)
      1'b0 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_2[31 : 0];
      default : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_2[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3_1)
      1'b0 : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_3[31 : 0];
      default : _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3 = execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_3[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_60)
      3'b000 : _zz_59 = _zz_45;
      3'b001 : _zz_59 = _zz_46;
      3'b010 : _zz_59 = _zz_47;
      3'b011 : _zz_59 = _zz_48;
      3'b100 : _zz_59 = _zz_49;
      3'b101 : _zz_59 = _zz_50;
      3'b110 : _zz_59 = _zz_51;
      default : _zz_59 = _zz_52;
    endcase
  end

  always @(*) begin
    case(_zz_62)
      3'b000 : _zz_61 = _zz_45;
      3'b001 : _zz_61 = _zz_46;
      3'b010 : _zz_61 = _zz_47;
      3'b011 : _zz_61 = _zz_48;
      3'b100 : _zz_61 = _zz_49;
      3'b101 : _zz_61 = _zz_50;
      3'b110 : _zz_61 = _zz_51;
      default : _zz_61 = _zz_52;
    endcase
  end

  always @(*) begin
    case(_zz_65)
      3'b000 : _zz_64 = 2'b00;
      3'b001 : _zz_64 = 2'b01;
      3'b010 : _zz_64 = 2'b01;
      3'b011 : _zz_64 = 2'b10;
      3'b100 : _zz_64 = 2'b01;
      3'b101 : _zz_64 = 2'b10;
      3'b110 : _zz_64 = 2'b10;
      default : _zz_64 = 2'b11;
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_lsu_ctrl_needFlushSel)
      2'b00 : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
      end
      2'b01 : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
      end
      2'b10 : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault;
      end
      default : begin
        _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address;
        _zz_LsuL1Plugin_logic_waysWrite_tag_fault = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault;
      end
    endcase
  end

  always @(*) begin
    case(LsuL1Plugin_logic_lsu_ctrl_targetWay)
      2'b00 : _zz_LsuL1Plugin_logic_writeback_push_payload_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
      2'b01 : _zz_LsuL1Plugin_logic_writeback_push_payload_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
      2'b10 : _zz_LsuL1Plugin_logic_writeback_push_payload_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address;
      default : _zz_LsuL1Plugin_logic_writeback_push_payload_address = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_1)
      2'b00 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_0;
      2'b01 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_1;
      2'b10 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_2;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted = LsuPlugin_logic_onCtrl_loadData_splitted_3;
    endcase
  end

  always @(*) begin
    case(_zz_LsuPlugin_logic_onCtrl_loadData_shifted_3)
      1'b0 : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_1;
      default : _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2 = LsuPlugin_logic_onCtrl_loadData_splitted_3;
    endcase
  end

  always @(*) begin
    case(LsuL1TileLinkPlugin_logic_down_a_payload_size)
      3'b000 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b000;
      3'b001 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b000;
      3'b010 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b000;
      3'b011 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b000;
      3'b100 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b001;
      3'b101 : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b011;
      default : _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last = 3'b111;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_0_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_0_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_0_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_1_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_1_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_1_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_2_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_2_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_2_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_3_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_3_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_3_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_4_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_4_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_4_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_5_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_5_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_5_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_6_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_6_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_6_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_7_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_7_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_7_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_8_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_8_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_8_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_9_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_9_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_9_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_10_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_10_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_10_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_11_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_11_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_11_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_12_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_12_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_12_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_PerformanceCounterPlugin_logic_events_sums_13_2)
      1'b0 : _zz_PerformanceCounterPlugin_logic_events_sums_13_1 = 1'b0;
      default : _zz_PerformanceCounterPlugin_logic_events_sums_13_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(CsrRamPlugin_logic_readLogic_sel)
      2'b00 : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = PerformanceCounterPlugin_logic_readPort_address;
      2'b01 : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = TrapPlugin_logic_harts_0_crsPorts_read_address;
      default : _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload = CsrRamPlugin_csrMapper_read_address;
    endcase
  end

  always @(*) begin
    case(_zz_WhiteboxerPlugin_logic_perf_candidatesCount_1)
      1'b0 : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 1'b0;
      default : _zz_WhiteboxerPlugin_logic_perf_candidatesCount = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount_1)
      1'b0 : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 1'b0;
      default : _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount = 1'b1;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : execute_ctrl2_up_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0)
      Input2Kind_RS : execute_ctrl2_up_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "RS   ";
      Input2Kind_IMM_I : execute_ctrl2_up_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "IMM_I";
      default : execute_ctrl2_up_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : execute_ctrl1_down_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0)
      Input2Kind_RS : execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "RS   ";
      Input2Kind_IMM_I : execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "IMM_I";
      default : execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0)
      Input2Kind_RS : execute_ctrl2_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "RS   ";
      Input2Kind_IMM_I : execute_ctrl2_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "IMM_I";
      default : execute_ctrl2_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_ECALL : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "ECALL     ";
      EnvPluginOp_EBREAK : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "SFENCE_VMA";
      EnvPluginOp_WFI : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "WFI       ";
      default : execute_ctrl2_down_early0_EnvPlugin_OP_lane0_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(FetchL1TileLinkPlugin_logic_down_a_payload_opcode)
      A_PUT_FULL_DATA : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : FetchL1TileLinkPlugin_logic_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(FetchL1TileLinkPlugin_logic_down_d_payload_opcode)
      D_ACCESS_ACK : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : FetchL1TileLinkPlugin_logic_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_ls_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_ls_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_access_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_access_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_onAddress0_flush_port_payload_op)
      LsuL1CmdOpcode_LSU : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "PREFETCH    ";
      default : LsuPlugin_logic_onAddress0_flush_port_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(LsuL1TileLinkPlugin_logic_down_a_payload_opcode)
      A_PUT_FULL_DATA : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : LsuL1TileLinkPlugin_logic_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(LsuL1TileLinkPlugin_logic_down_d_payload_opcode)
      D_ACCESS_ACK : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : LsuL1TileLinkPlugin_logic_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode)
      A_PUT_FULL_DATA : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode)
      D_ACCESS_ACK : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "RELEASE_ACK    ";
      default : LsuTileLinkPlugin_logic_bridge_down_d_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode)
      A_PUT_FULL_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2)
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "XOR_1";
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "OR_1 ";
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "AND_1";
      IntAluPlugin_AluBitwiseCtrlEnum_ZERO : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "ZERO ";
      default : _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2)
      BranchPlugin_BranchCtrlEnum_B : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "B   ";
      BranchPlugin_BranchCtrlEnum_JAL : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "JAL ";
      BranchPlugin_BranchCtrlEnum_JALR : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "JALR";
      default : _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0)
      Input2Kind_RS : _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "RS   ";
      Input2Kind_IMM_I : _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "IMM_I";
      default : _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_1)
      Input2Kind_RS : _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_1_string = "RS   ";
      Input2Kind_IMM_I : _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_1_string = "IMM_I";
      default : _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_2)
      Input2Kind_RS : _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_2_string = "RS   ";
      Input2Kind_IMM_I : _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_2_string = "IMM_I";
      default : _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1)
      EnvPluginOp_ECALL : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "WFI       ";
      default : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2)
      EnvPluginOp_ECALL : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "WFI       ";
      default : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3)
      EnvPluginOp_ECALL : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "ECALL     ";
      EnvPluginOp_EBREAK : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "EBREAK    ";
      EnvPluginOp_PRIV_RET : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "PRIV_RET  ";
      EnvPluginOp_FENCE_I : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "FENCE_I   ";
      EnvPluginOp_SFENCE_VMA : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "SFENCE_VMA";
      EnvPluginOp_WFI : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "WFI       ";
      default : _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3_string = "??????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_IDLE : LsuPlugin_logic_flusher_stateReg_string = "IDLE      ";
      LsuPlugin_logic_flusher_CMD : LsuPlugin_logic_flusher_stateReg_string = "CMD       ";
      LsuPlugin_logic_flusher_COMPLETION : LsuPlugin_logic_flusher_stateReg_string = "COMPLETION";
      default : LsuPlugin_logic_flusher_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(LsuPlugin_logic_flusher_stateNext)
      LsuPlugin_logic_flusher_IDLE : LsuPlugin_logic_flusher_stateNext_string = "IDLE      ";
      LsuPlugin_logic_flusher_CMD : LsuPlugin_logic_flusher_stateNext_string = "CMD       ";
      LsuPlugin_logic_flusher_COMPLETION : LsuPlugin_logic_flusher_stateNext_string = "COMPLETION";
      default : LsuPlugin_logic_flusher_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RESET : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "RESET      ";
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "RUNNING    ";
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "PROCESS_1  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_TVAL  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_TVEC  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "TRAP_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "XRET_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "XRET_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "ATS_RSP    ";
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "JUMP       ";
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "LSU_FLUSH  ";
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "FETCH_FLUSH";
      default : TrapPlugin_logic_harts_0_trap_fsm_stateReg_string = "???????????";
    endcase
  end
  always @(*) begin
    case(TrapPlugin_logic_harts_0_trap_fsm_stateNext)
      TrapPlugin_logic_harts_0_trap_fsm_RESET : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "RESET      ";
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "RUNNING    ";
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "PROCESS_1  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_TVAL  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_TVEC  ";
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "TRAP_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "XRET_EPC   ";
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "XRET_APPLY ";
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "ATS_RSP    ";
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "JUMP       ";
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "LSU_FLUSH  ";
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "FETCH_FLUSH";
      default : TrapPlugin_logic_harts_0_trap_fsm_stateNext_string = "???????????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_BOOT : MmuPlugin_logic_refill_stateReg_string = "BOOT ";
      MmuPlugin_logic_refill_IDLE : MmuPlugin_logic_refill_stateReg_string = "IDLE ";
      MmuPlugin_logic_refill_CMD_0 : MmuPlugin_logic_refill_stateReg_string = "CMD_0";
      MmuPlugin_logic_refill_CMD_1 : MmuPlugin_logic_refill_stateReg_string = "CMD_1";
      MmuPlugin_logic_refill_RSP_0 : MmuPlugin_logic_refill_stateReg_string = "RSP_0";
      MmuPlugin_logic_refill_RSP_1 : MmuPlugin_logic_refill_stateReg_string = "RSP_1";
      default : MmuPlugin_logic_refill_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(MmuPlugin_logic_refill_stateNext)
      MmuPlugin_logic_refill_BOOT : MmuPlugin_logic_refill_stateNext_string = "BOOT ";
      MmuPlugin_logic_refill_IDLE : MmuPlugin_logic_refill_stateNext_string = "IDLE ";
      MmuPlugin_logic_refill_CMD_0 : MmuPlugin_logic_refill_stateNext_string = "CMD_0";
      MmuPlugin_logic_refill_CMD_1 : MmuPlugin_logic_refill_stateNext_string = "CMD_1";
      MmuPlugin_logic_refill_RSP_0 : MmuPlugin_logic_refill_stateNext_string = "RSP_0";
      MmuPlugin_logic_refill_RSP_1 : MmuPlugin_logic_refill_stateNext_string = "RSP_1";
      default : MmuPlugin_logic_refill_stateNext_string = "?????";
    endcase
  end
  always @(*) begin
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_BOOT : PerformanceCounterPlugin_logic_fsm_stateReg_string = "BOOT     ";
      PerformanceCounterPlugin_logic_fsm_IDLE : PerformanceCounterPlugin_logic_fsm_stateReg_string = "IDLE     ";
      PerformanceCounterPlugin_logic_fsm_READ_LOW : PerformanceCounterPlugin_logic_fsm_stateReg_string = "READ_LOW ";
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : PerformanceCounterPlugin_logic_fsm_stateReg_string = "CALC_LOW ";
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : PerformanceCounterPlugin_logic_fsm_stateReg_string = "READ_HIGH";
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : PerformanceCounterPlugin_logic_fsm_stateReg_string = "CALC_HIGH";
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : PerformanceCounterPlugin_logic_fsm_stateReg_string = "CSR_WRITE";
      default : PerformanceCounterPlugin_logic_fsm_stateReg_string = "?????????";
    endcase
  end
  always @(*) begin
    case(PerformanceCounterPlugin_logic_fsm_stateNext)
      PerformanceCounterPlugin_logic_fsm_BOOT : PerformanceCounterPlugin_logic_fsm_stateNext_string = "BOOT     ";
      PerformanceCounterPlugin_logic_fsm_IDLE : PerformanceCounterPlugin_logic_fsm_stateNext_string = "IDLE     ";
      PerformanceCounterPlugin_logic_fsm_READ_LOW : PerformanceCounterPlugin_logic_fsm_stateNext_string = "READ_LOW ";
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : PerformanceCounterPlugin_logic_fsm_stateNext_string = "CALC_LOW ";
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : PerformanceCounterPlugin_logic_fsm_stateNext_string = "READ_HIGH";
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : PerformanceCounterPlugin_logic_fsm_stateNext_string = "CALC_HIGH";
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : PerformanceCounterPlugin_logic_fsm_stateNext_string = "CSR_WRITE";
      default : PerformanceCounterPlugin_logic_fsm_stateNext_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_IDLE : CsrAccessPlugin_logic_fsm_stateReg_string = "IDLE      ";
      CsrAccessPlugin_logic_fsm_READ : CsrAccessPlugin_logic_fsm_stateReg_string = "READ      ";
      CsrAccessPlugin_logic_fsm_WRITE : CsrAccessPlugin_logic_fsm_stateReg_string = "WRITE     ";
      CsrAccessPlugin_logic_fsm_COMPLETION : CsrAccessPlugin_logic_fsm_stateReg_string = "COMPLETION";
      default : CsrAccessPlugin_logic_fsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(CsrAccessPlugin_logic_fsm_stateNext)
      CsrAccessPlugin_logic_fsm_IDLE : CsrAccessPlugin_logic_fsm_stateNext_string = "IDLE      ";
      CsrAccessPlugin_logic_fsm_READ : CsrAccessPlugin_logic_fsm_stateNext_string = "READ      ";
      CsrAccessPlugin_logic_fsm_WRITE : CsrAccessPlugin_logic_fsm_stateNext_string = "WRITE     ";
      CsrAccessPlugin_logic_fsm_COMPLETION : CsrAccessPlugin_logic_fsm_stateNext_string = "COMPLETION";
      default : CsrAccessPlugin_logic_fsm_stateNext_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    BtbPlugin_logic_ras_ptr_pop_aheadValue = BtbPlugin_logic_ras_ptr_pop;
    BtbPlugin_logic_ras_ptr_pop_aheadValue = (_zz_BtbPlugin_logic_ras_ptr_pop_aheadValue - _zz_BtbPlugin_logic_ras_ptr_pop_aheadValue_3);
  end

  assign execute_ctrl4_down_RD_ENABLE_lane0 = execute_ctrl4_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl4_RD_ENABLE_lane0_bypass = execute_ctrl4_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_4) begin
      execute_ctrl4_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl4_down_LANE_SEL_lane0 = execute_ctrl4_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl4_LANE_SEL_lane0_bypass = execute_ctrl4_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_4) begin
      execute_ctrl4_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_RD_ENABLE_lane0 = execute_ctrl3_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl3_RD_ENABLE_lane0_bypass = execute_ctrl3_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_3) begin
      execute_ctrl3_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_LANE_SEL_lane0 = execute_ctrl3_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl3_LANE_SEL_lane0_bypass = execute_ctrl3_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_3) begin
      execute_ctrl3_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl2_down_RD_ENABLE_lane0 = execute_ctrl2_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl2_RD_ENABLE_lane0_bypass = execute_ctrl2_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_2) begin
      execute_ctrl2_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl2_down_LANE_SEL_lane0 = execute_ctrl2_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl2_LANE_SEL_lane0_bypass = execute_ctrl2_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_2) begin
      execute_ctrl2_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl1_down_RD_ENABLE_lane0 = execute_ctrl1_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl1_RD_ENABLE_lane0_bypass = execute_ctrl1_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306_1) begin
      execute_ctrl1_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl1_down_LANE_SEL_lane0 = execute_ctrl1_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl1_LANE_SEL_lane0_bypass = execute_ctrl1_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306_1) begin
      execute_ctrl1_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl0_down_RD_ENABLE_lane0 = execute_ctrl0_RD_ENABLE_lane0_bypass;
  always @(*) begin
    execute_ctrl0_RD_ENABLE_lane0_bypass = execute_ctrl0_up_RD_ENABLE_lane0;
    if(when_ExecuteLanePlugin_l306) begin
      execute_ctrl0_RD_ENABLE_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl0_down_LANE_SEL_lane0 = execute_ctrl0_LANE_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl0_LANE_SEL_lane0_bypass = execute_ctrl0_up_LANE_SEL_lane0;
    if(when_ExecuteLanePlugin_l306) begin
      execute_ctrl0_LANE_SEL_lane0_bypass = 1'b0;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(CsrRamPlugin_logic_writeLogic_port_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    PcPlugin_logic_harts_0_aggregator_fault_1 = PcPlugin_logic_harts_0_aggregator_fault;
    if(when_PcPlugin_l80) begin
      PcPlugin_logic_harts_0_aggregator_fault_1 = _zz_PcPlugin_logic_harts_0_aggregator_fault_1_1[0];
    end
  end

  always @(*) begin
    PcPlugin_logic_harts_0_aggregator_target_1 = PcPlugin_logic_harts_0_aggregator_target;
    if(when_PcPlugin_l80) begin
      PcPlugin_logic_harts_0_aggregator_target_1 = (_zz_PcPlugin_logic_harts_0_aggregator_fault_1 ? BtbPlugin_logic_pcPort_payload_pc : 32'h0);
    end
  end

  assign execute_ctrl4_down_COMMIT_lane0 = execute_ctrl4_COMMIT_lane0_bypass;
  always @(*) begin
    execute_ctrl4_COMMIT_lane0_bypass = execute_ctrl4_up_COMMIT_lane0;
    if(when_LsuPlugin_l861) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        execute_ctrl4_COMMIT_lane0_bypass = 1'b0;
      end
    end
  end

  assign execute_ctrl4_down_TRAP_lane0 = execute_ctrl4_TRAP_lane0_bypass;
  always @(*) begin
    execute_ctrl4_TRAP_lane0_bypass = execute_ctrl4_up_TRAP_lane0;
    if(when_LsuPlugin_l861) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        execute_ctrl4_TRAP_lane0_bypass = 1'b1;
      end
    end
  end

  assign execute_ctrl4_down_LsuL1_SEL_lane0 = execute_ctrl4_LsuL1_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl4_LsuL1_SEL_lane0_bypass = execute_ctrl4_up_LsuL1_SEL_lane0;
    if(when_LsuPlugin_l546_1) begin
      execute_ctrl4_LsuL1_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_LsuL1_SEL_lane0 = execute_ctrl3_LsuL1_SEL_lane0_bypass;
  always @(*) begin
    execute_ctrl3_LsuL1_SEL_lane0_bypass = execute_ctrl3_up_LsuL1_SEL_lane0;
    if(when_LsuPlugin_l546) begin
      execute_ctrl3_LsuL1_SEL_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0 = execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_1 = execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_1;
  assign execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty = execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty;
  always @(*) begin
    _zz_3 = 1'b0;
    if(LsuL1Plugin_logic_writeback_read_slotReadLast_valid) begin
      _zz_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_4 = 1'b0;
    if(LsuL1Plugin_logic_shared_write_valid) begin
      _zz_4 = 1'b1;
    end
  end

  assign decode_ctrls_1_down_LANE_SEL_0 = decode_ctrls_1_LANE_SEL_0_bypass;
  always @(*) begin
    decode_ctrls_1_LANE_SEL_0_bypass = decode_ctrls_1_up_LANE_SEL_0;
    if(decode_logic_flushes_1_onLanes_0_doIt) begin
      decode_ctrls_1_LANE_SEL_0_bypass = 1'b0;
    end
  end

  assign decode_ctrls_0_down_LANE_SEL_0 = decode_ctrls_0_LANE_SEL_0_bypass;
  always @(*) begin
    decode_ctrls_0_LANE_SEL_0_bypass = decode_ctrls_0_up_LANE_SEL_0;
    if(decode_logic_flushes_0_onLanes_0_doIt) begin
      decode_ctrls_0_LANE_SEL_0_bypass = 1'b0;
    end
  end

  assign execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass;
  assign decode_ctrls_1_down_TRAP_0 = decode_ctrls_1_TRAP_0_bypass;
  always @(*) begin
    decode_ctrls_1_TRAP_0_bypass = decode_ctrls_1_up_TRAP_0;
    if(when_DecoderPlugin_l229) begin
      decode_ctrls_1_TRAP_0_bypass = 1'b1;
    end
  end

  assign execute_ctrl4_down_COMPLETED_lane0 = execute_ctrl4_COMPLETED_lane0_bypass;
  assign execute_ctrl3_down_COMPLETED_lane0 = execute_ctrl3_COMPLETED_lane0_bypass;
  assign execute_ctrl2_down_COMPLETED_lane0 = execute_ctrl2_COMPLETED_lane0_bypass;
  assign execute_ctrl3_down_COMMIT_lane0 = execute_ctrl3_COMMIT_lane0_bypass;
  always @(*) begin
    execute_ctrl3_COMMIT_lane0_bypass = execute_ctrl3_up_COMMIT_lane0;
    if(when_BranchPlugin_l251) begin
      execute_ctrl3_COMMIT_lane0_bypass = 1'b0;
    end
  end

  assign execute_ctrl3_down_TRAP_lane0 = execute_ctrl3_TRAP_lane0_bypass;
  always @(*) begin
    execute_ctrl3_TRAP_lane0_bypass = execute_ctrl3_up_TRAP_lane0;
    if(when_BranchPlugin_l251) begin
      execute_ctrl3_TRAP_lane0_bypass = 1'b1;
    end
  end

  always @(*) begin
    early0_BranchPlugin_logic_jumpLogic_history_shifter_1 = early0_BranchPlugin_logic_jumpLogic_history_shifter;
    if(when_BranchPlugin_l218) begin
      early0_BranchPlugin_logic_jumpLogic_history_shifter_1 = _zz_early0_BranchPlugin_logic_jumpLogic_history_shifter_1[11 : 0];
    end
  end

  assign execute_ctrl2_down_COMMIT_lane0 = execute_ctrl2_COMMIT_lane0_bypass;
  always @(*) begin
    execute_ctrl2_COMMIT_lane0_bypass = execute_ctrl2_up_COMMIT_lane0;
    if(when_EnvPlugin_l119) begin
      if(when_EnvPlugin_l123) begin
        execute_ctrl2_COMMIT_lane0_bypass = 1'b0;
      end
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              execute_ctrl2_COMMIT_lane0_bypass = 1'b0;
            end
          end
        end
      end
    endcase
  end

  assign execute_ctrl2_down_TRAP_lane0 = execute_ctrl2_TRAP_lane0_bypass;
  always @(*) begin
    execute_ctrl2_TRAP_lane0_bypass = execute_ctrl2_up_TRAP_lane0;
    if(when_EnvPlugin_l119) begin
      execute_ctrl2_TRAP_lane0_bypass = 1'b1;
    end
    if(CsrAccessPlugin_logic_fsm_inject_flushReg) begin
      execute_ctrl2_TRAP_lane0_bypass = 1'b1;
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              execute_ctrl2_TRAP_lane0_bypass = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                execute_ctrl2_TRAP_lane0_bypass = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    _zz_wr_en = 1'b0;
    if(BtbPlugin_logic_ras_write_valid) begin
      _zz_wr_en = 1'b1;
    end
  end

  always @(*) begin
    _zz_5 = 1'b0;
    if(GSharePlugin_logic_mem_write_valid) begin
      _zz_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217 = 1'b0;
    if(when_FetchL1Plugin_l216) begin
      _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217 = 1'b1;
    end
  end

  always @(*) begin
    _zz_6 = 1'b0;
    if(FetchL1Plugin_logic_plru_write_valid) begin
      _zz_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_7 = 1'b0;
    if(FetchL1Plugin_logic_banks_3_write_valid) begin
      _zz_7 = 1'b1;
    end
  end

  always @(*) begin
    _zz_8 = 1'b0;
    if(FetchL1Plugin_logic_banks_2_write_valid) begin
      _zz_8 = 1'b1;
    end
  end

  always @(*) begin
    _zz_9 = 1'b0;
    if(FetchL1Plugin_logic_banks_1_write_valid) begin
      _zz_9 = 1'b1;
    end
  end

  always @(*) begin
    _zz_10 = 1'b0;
    if(FetchL1Plugin_logic_banks_0_write_valid) begin
      _zz_10 = 1'b1;
    end
  end

  assign AlignerPlugin_api_singleFetch = 1'b0;
  assign AlignerPlugin_api_haltIt = 1'b0;
  always @(*) begin
    DispatchPlugin_api_haltDispatch = 1'b0;
    if(LsuPlugin_logic_onCtrl_hartRegulation_valid) begin
      DispatchPlugin_api_haltDispatch = 1'b1;
    end
  end

  always @(*) begin
    CsrRamPlugin_api_holdRead = 1'b0;
    if(PerformanceCounterPlugin_logic_csrRead_requested) begin
      if(when_PerformanceCounterPlugin_l342) begin
        CsrRamPlugin_api_holdRead = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrRamPlugin_api_holdWrite = 1'b0;
    if(PerformanceCounterPlugin_logic_fsm_holdCsrWrite) begin
      CsrRamPlugin_api_holdWrite = 1'b1;
    end
  end

  always @(*) begin
    TrapPlugin_api_harts_0_redo = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
              TrapPlugin_api_harts_0_redo = 1'b1;
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
        if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid) begin
          TrapPlugin_api_harts_0_redo = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_api_harts_0_askWake = 1'b0;
    if(when_TrapPlugin_l226) begin
      TrapPlugin_api_harts_0_askWake = 1'b1;
    end
  end

  always @(*) begin
    TrapPlugin_api_harts_0_rvTrap = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_api_harts_0_rvTrap = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0)
      IntAluPlugin_AluBitwiseCtrlEnum_AND_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 & execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_OR_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 | execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      IntAluPlugin_AluBitwiseCtrlEnum_XOR_1 : begin
        early0_IntAluPlugin_logic_alu_bitwise = (execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 ^ execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
      end
      default : begin
        early0_IntAluPlugin_logic_alu_bitwise = 32'h0;
      end
    endcase
  end

  assign early0_IntAluPlugin_logic_alu_result = (_zz_early0_IntAluPlugin_logic_alu_result | _zz_early0_IntAluPlugin_logic_alu_result_2);
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0 = early0_IntAluPlugin_logic_alu_result;
  assign early0_IntAluPlugin_logic_wb_valid = execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0;
  assign early0_IntAluPlugin_logic_wb_payload = execute_ctrl2_down_early0_IntAluPlugin_ALU_RESULT_lane0;
  assign early0_BarrelShifterPlugin_logic_shift_amplitude = _zz_early0_BarrelShifterPlugin_logic_shift_amplitude;
  assign early0_BarrelShifterPlugin_logic_shift_reversed = (execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_early0_BarrelShifterPlugin_logic_shift_reversed : execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0);
  assign early0_BarrelShifterPlugin_logic_shift_shifted = _zz_early0_BarrelShifterPlugin_logic_shift_shifted[31:0];
  assign early0_BarrelShifterPlugin_logic_shift_patched = (execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 ? _zz_early0_BarrelShifterPlugin_logic_shift_patched : early0_BarrelShifterPlugin_logic_shift_shifted);
  assign execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0 = early0_BarrelShifterPlugin_logic_shift_patched;
  assign early0_BarrelShifterPlugin_logic_wb_valid = execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0;
  assign early0_BarrelShifterPlugin_logic_wb_payload = execute_ctrl2_down_early0_BarrelShifterPlugin_SHIFT_RESULT_lane0;
  assign CfuPlugin_logic_onFork_schedule = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CfuPlugin_logic_CFU_ENABLE_lane0);
  assign CfuPlugin_logic_onFork_hold = 1'b0;
  assign CfuPlugin_logic_bus_cmd_fire = (CfuPlugin_logic_bus_cmd_valid && CfuPlugin_logic_bus_cmd_ready);
  assign when_CfuPlugin_l147 = (! execute_freeze_valid);
  assign execute_ctrl2_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0 = ((CfuPlugin_logic_onFork_schedule || CfuPlugin_logic_onFork_hold) || CfuPlugin_logic_onFork_fired);
  assign CfuPlugin_logic_bus_cmd_valid = ((CfuPlugin_logic_onFork_schedule || CfuPlugin_logic_onFork_hold) && (! CfuPlugin_logic_onFork_fired));
  assign CfuPlugin_logic_onFork_freezeIt = (CfuPlugin_logic_bus_cmd_valid && (! CfuPlugin_logic_bus_cmd_ready));
  always @(*) begin
    LsuPlugin_logic_events_waiting = 1'b0;
    if(LsuPlugin_logic_onCtrl_hartRegulation_valid) begin
      LsuPlugin_logic_events_waiting = 1'b1;
    end
  end

  always @(*) begin
    LsuL1_ackUnlock = 1'b0;
    if(LsuPlugin_logic_onCtrl_io_cmdSent) begin
      LsuL1_ackUnlock = 1'b1;
    end
  end

  assign execute_ctrl2_down_MUL_SRC1_lane0 = _zz_execute_ctrl2_down_MUL_SRC1_lane0;
  assign execute_ctrl2_down_MUL_SRC2_lane0 = _zz_execute_ctrl2_down_MUL_SRC2_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = (execute_ctrl2_down_MUL_SRC1_lane0[16 : 0] * execute_ctrl2_down_MUL_SRC2_lane0[16 : 0]);
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = _zz_execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[33 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0[33 : 0];
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[60 : 34] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0[26 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_1[60 : 17] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0[43 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2 = 61'h0;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_2[60 : 17] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0[43 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0[29 : 27];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_1[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0[46 : 44];
  end

  always @(*) begin
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2 = 3'b000;
    _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_2[2 : 0] = execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0[46 : 44];
  end

  assign execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_3 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0_6);
  assign execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = (_zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_3 + _zz_execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0_6);
  always @(*) begin
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 = 66'h0;
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[62 : 0] = execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0[62 : 0];
  end

  always @(*) begin
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1 = 66'h0;
    _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1[65 : 61] = execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0[4 : 0];
  end

  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 = (_zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0 + _zz_execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0_1);
  assign early0_MulPlugin_logic_formatBus_valid = execute_ctrl4_down_early0_MulPlugin_SEL_lane0;
  assign early0_MulPlugin_logic_formatBus_payload = (execute_ctrl4_down_MulPlugin_HIGH_lane0 ? execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[63 : 32] : execute_ctrl4_down_early0_MulPlugin_logic_steps_1_adders_0_lane0[31 : 0]);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0 = execute_ctrl2_up_integer_RS1_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0 = execute_ctrl2_up_integer_RS2_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 = (execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 && execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0[31]);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 = (execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 && execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0[31]);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0 = ((execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 ? (~ execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0) : execute_ctrl2_down_RsUnsignedPlugin_RS1_FORMATED_lane0) + _zz_execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0);
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0 = ((execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 ? (~ execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0) : execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0) + _zz_execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0);
  assign early0_DivPlugin_logic_processing_div_io_cmd_fire = (early0_DivPlugin_logic_processing_div_io_cmd_valid && early0_DivPlugin_logic_processing_div_io_cmd_ready);
  assign early0_DivPlugin_logic_processing_request = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_early0_DivPlugin_SEL_lane0);
  assign early0_DivPlugin_logic_processing_a = execute_ctrl2_down_RsUnsignedPlugin_RS1_UNSIGNED_lane0;
  assign early0_DivPlugin_logic_processing_b = execute_ctrl2_down_RsUnsignedPlugin_RS2_UNSIGNED_lane0;
  assign early0_DivPlugin_logic_processing_div_io_cmd_valid = (early0_DivPlugin_logic_processing_request && (! early0_DivPlugin_logic_processing_cmdSent));
  assign early0_DivPlugin_logic_processing_freeze = ((early0_DivPlugin_logic_processing_request && (! early0_DivPlugin_logic_processing_div_io_rsp_valid)) && (! early0_DivPlugin_logic_processing_unscheduleRequest));
  assign early0_DivPlugin_logic_processing_selected = (execute_ctrl2_down_DivPlugin_REM_lane0 ? early0_DivPlugin_logic_processing_div_io_rsp_payload_remain : early0_DivPlugin_logic_processing_div_io_rsp_payload_result);
  assign _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0 = early0_DivPlugin_logic_processing_selected;
  assign execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0 = _zz_execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0_1;
  assign early0_DivPlugin_logic_formatBus_valid = execute_ctrl3_down_early0_DivPlugin_SEL_lane0;
  assign early0_DivPlugin_logic_formatBus_payload = execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0;
  assign WhiteboxerPlugin_logic_fetch_fire = fetch_logic_ctrls_0_down_isFiring;
  assign PrivilegedPlugin_api_harts_0_allowInterrupts = 1'b1;
  assign PrivilegedPlugin_api_harts_0_allowException = 1'b1;
  assign PrivilegedPlugin_api_harts_0_allowEbreakException = 1'b1;
  assign PrivilegedPlugin_api_harts_0_fpuEnable = 1'b0;
  always @(*) begin
    CsrAccessPlugin_bus_decode_exception = 1'b0;
    if(when_PrivilegedPlugin_l689) begin
      CsrAccessPlugin_bus_decode_exception = 1'b1;
    end
    if(when_CsrAccessPlugin_l155) begin
      if(when_MmuPlugin_l221) begin
        CsrAccessPlugin_bus_decode_exception = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l155_2) begin
      if(when_PerformanceCounterPlugin_l327) begin
        if(when_PerformanceCounterPlugin_l328) begin
          CsrAccessPlugin_bus_decode_exception = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_decode_trap = 1'b0;
    if(when_CsrAccessPlugin_l155) begin
      if(!when_MmuPlugin_l221) begin
        CsrAccessPlugin_bus_decode_trap = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l155_1) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trap = 1'b1;
      end
    end
    if(when_CsrAccessPlugin_l155_3) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trap = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_decode_trapCode = 4'bxxxx;
    if(when_CsrAccessPlugin_l155) begin
      if(!when_MmuPlugin_l221) begin
        CsrAccessPlugin_bus_decode_trapCode = 4'b0110;
      end
    end
    if(when_CsrAccessPlugin_l155_1) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trapCode = 4'b0101;
      end
    end
    if(when_CsrAccessPlugin_l155_3) begin
      if(CsrAccessPlugin_bus_decode_write) begin
        CsrAccessPlugin_bus_decode_trapCode = 4'b0101;
      end
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_read_halt = 1'b0;
    if(when_CsrRamPlugin_l85) begin
      CsrAccessPlugin_bus_read_halt = 1'b1;
    end
  end

  always @(*) begin
    CsrAccessPlugin_bus_write_halt = 1'b0;
    if(when_CsrRamPlugin_l96) begin
      CsrAccessPlugin_bus_write_halt = 1'b1;
    end
    if(when_CsrAccessPlugin_l343_3) begin
      if(when_PerformanceCounterPlugin_l357) begin
        if(when_PerformanceCounterPlugin_l359) begin
          CsrAccessPlugin_bus_write_halt = 1'b1;
        end
      end
    end
  end

  assign FetchL1Plugin_logic_banks_0_read_rsp = FetchL1Plugin_logic_banks_0_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_0 = FetchL1Plugin_logic_banks_0_read_rsp;
  assign FetchL1Plugin_logic_banks_1_read_rsp = FetchL1Plugin_logic_banks_1_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_1 = FetchL1Plugin_logic_banks_1_read_rsp;
  assign FetchL1Plugin_logic_banks_2_read_rsp = FetchL1Plugin_logic_banks_2_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_2 = FetchL1Plugin_logic_banks_2_read_rsp;
  assign FetchL1Plugin_logic_banks_3_read_rsp = FetchL1Plugin_logic_banks_3_mem_spinal_port1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_WORDS_3 = FetchL1Plugin_logic_banks_3_read_rsp;
  always @(*) begin
    FetchL1Plugin_logic_waysWrite_mask = 4'b0000;
    if(when_FetchL1Plugin_l204) begin
      FetchL1Plugin_logic_waysWrite_mask = 4'b1111;
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      if(when_FetchL1Plugin_l304) begin
        FetchL1Plugin_logic_waysWrite_mask[FetchL1Plugin_logic_refill_onRsp_wayToAllocate] = 1'b1;
      end
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_address = 6'bxxxxxx;
    if(when_FetchL1Plugin_l204) begin
      FetchL1Plugin_logic_waysWrite_address = FetchL1Plugin_logic_invalidate_counter[5:0];
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_address = FetchL1Plugin_logic_refill_onRsp_address[11 : 6];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_loaded = 1'bx;
    if(when_FetchL1Plugin_l204) begin
      FetchL1Plugin_logic_waysWrite_tag_loaded = 1'b0;
    end
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_error = 1'bx;
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_error = (FetchL1Plugin_logic_bus_rsp_valid && FetchL1Plugin_logic_bus_rsp_payload_error);
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(FetchL1Plugin_logic_invalidate_done) begin
      FetchL1Plugin_logic_waysWrite_tag_address = FetchL1Plugin_logic_refill_onRsp_address[31 : 12];
    end
  end

  assign _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded = FetchL1Plugin_logic_ways_0_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_0_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_0_read_rsp_error = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_0_read_rsp_address = _zz_FetchL1Plugin_logic_ways_0_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded = FetchL1Plugin_logic_ways_0_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error = FetchL1Plugin_logic_ways_0_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address = FetchL1Plugin_logic_ways_0_read_rsp_address;
  assign _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded = FetchL1Plugin_logic_ways_1_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_1_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_1_read_rsp_error = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_1_read_rsp_address = _zz_FetchL1Plugin_logic_ways_1_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded = FetchL1Plugin_logic_ways_1_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error = FetchL1Plugin_logic_ways_1_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address = FetchL1Plugin_logic_ways_1_read_rsp_address;
  assign _zz_FetchL1Plugin_logic_ways_2_read_rsp_loaded = FetchL1Plugin_logic_ways_2_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_2_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_2_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_2_read_rsp_error = _zz_FetchL1Plugin_logic_ways_2_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_2_read_rsp_address = _zz_FetchL1Plugin_logic_ways_2_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_loaded = FetchL1Plugin_logic_ways_2_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_error = FetchL1Plugin_logic_ways_2_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_address = FetchL1Plugin_logic_ways_2_read_rsp_address;
  assign _zz_FetchL1Plugin_logic_ways_3_read_rsp_loaded = FetchL1Plugin_logic_ways_3_mem_spinal_port1;
  assign FetchL1Plugin_logic_ways_3_read_rsp_loaded = _zz_FetchL1Plugin_logic_ways_3_read_rsp_loaded[0];
  assign FetchL1Plugin_logic_ways_3_read_rsp_error = _zz_FetchL1Plugin_logic_ways_3_read_rsp_loaded[1];
  assign FetchL1Plugin_logic_ways_3_read_rsp_address = _zz_FetchL1Plugin_logic_ways_3_read_rsp_loaded[21 : 2];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_loaded = FetchL1Plugin_logic_ways_3_read_rsp_loaded;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_error = FetchL1Plugin_logic_ways_3_read_rsp_error;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_address = FetchL1Plugin_logic_ways_3_read_rsp_address;
  assign _zz_FetchL1Plugin_logic_plru_read_rsp_0 = FetchL1Plugin_logic_plru_mem_spinal_port1;
  assign FetchL1Plugin_logic_plru_read_rsp_0 = _zz_FetchL1Plugin_logic_plru_read_rsp_0[0 : 0];
  assign FetchL1Plugin_logic_plru_read_rsp_1 = _zz_FetchL1Plugin_logic_plru_read_rsp_0[2 : 1];
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0 = FetchL1Plugin_logic_plru_read_rsp_0;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_1 = FetchL1Plugin_logic_plru_read_rsp_1;
  assign FetchL1Plugin_logic_invalidate_cmd_valid = (|TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid);
  always @(*) begin
    FetchL1Plugin_logic_invalidate_canStart = 1'b1;
    if(when_FetchL1Plugin_l268) begin
      FetchL1Plugin_logic_invalidate_canStart = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_invalidate_counterIncr = (FetchL1Plugin_logic_invalidate_counter + 7'h01);
  assign FetchL1Plugin_logic_invalidate_done = FetchL1Plugin_logic_invalidate_counter[6];
  assign FetchL1Plugin_logic_invalidate_last = FetchL1Plugin_logic_invalidate_counterIncr[6];
  assign when_FetchL1Plugin_l204 = (! FetchL1Plugin_logic_invalidate_done);
  assign when_FetchL1Plugin_l211 = ((FetchL1Plugin_logic_invalidate_done && FetchL1Plugin_logic_invalidate_cmd_valid) && FetchL1Plugin_logic_invalidate_canStart);
  always @(*) begin
    TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready = 1'b0;
    if(when_FetchL1Plugin_l216) begin
      if(FetchL1Plugin_logic_invalidate_last) begin
        TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready = 1'b1;
      end
    end
  end

  assign when_FetchL1Plugin_l216 = (! FetchL1Plugin_logic_invalidate_done);
  assign fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217 = _zz_fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217;
  assign FetchL1Plugin_logic_refill_slots_0_askCmd = (FetchL1Plugin_logic_refill_slots_0_valid && (! FetchL1Plugin_logic_refill_slots_0_cmdSent));
  assign FetchL1Plugin_logic_refill_hazard = (|(FetchL1Plugin_logic_refill_slots_0_valid && (FetchL1Plugin_logic_refill_slots_0_address[11 : 6] == FetchL1Plugin_logic_refill_start_address[11 : 6])));
  assign when_FetchL1Plugin_l255 = ((FetchL1Plugin_logic_refill_start_valid && FetchL1Plugin_logic_invalidate_done) && (! FetchL1Plugin_logic_refill_hazard));
  assign when_FetchL1Plugin_l268 = ((|FetchL1Plugin_logic_refill_slots_0_valid) || FetchL1Plugin_logic_refill_start_valid);
  assign FetchL1Plugin_logic_refill_onCmd_propoedOh = (FetchL1Plugin_logic_refill_slots_0_askCmd && 1'b1);
  assign when_FetchL1Plugin_l276 = (! FetchL1Plugin_logic_refill_onCmd_locked);
  assign FetchL1Plugin_logic_refill_onCmd_oh = (FetchL1Plugin_logic_refill_onCmd_locked ? FetchL1Plugin_logic_refill_onCmd_lockedOh : FetchL1Plugin_logic_refill_onCmd_propoedOh);
  assign FetchL1Plugin_logic_bus_cmd_valid = (|FetchL1Plugin_logic_refill_onCmd_oh);
  assign FetchL1Plugin_logic_bus_cmd_payload_address = {FetchL1Plugin_logic_refill_slots_0_address[31 : 6],6'h0};
  assign FetchL1Plugin_logic_bus_cmd_payload_io = FetchL1Plugin_logic_refill_slots_0_isIo;
  assign FetchL1Plugin_logic_refill_onRsp_holdHarts = ((|FetchL1Plugin_logic_waysWrite_mask) || (|((FetchL1Plugin_logic_refill_slots_0_valid && (FetchL1Plugin_logic_refill_slots_0_address[11 : 6] == fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6])) && (! (1'b1 && (fetch_logic_ctrls_0_down_Fetch_WORD_PC[5 : 3] < FetchL1Plugin_logic_refill_onRsp_wordIndex))))));
  assign fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l297 = FetchL1Plugin_logic_refill_onRsp_holdHarts;
  assign FetchL1Plugin_logic_bus_rsp_fire = (FetchL1Plugin_logic_bus_rsp_valid && FetchL1Plugin_logic_bus_rsp_ready);
  assign FetchL1Plugin_logic_refill_onRsp_wayToAllocate = FetchL1Plugin_logic_refill_slots_0_wayToAllocate;
  assign FetchL1Plugin_logic_refill_onRsp_address = FetchL1Plugin_logic_refill_slots_0_address;
  assign when_FetchL1Plugin_l304 = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_firstCycle || FetchL1Plugin_logic_bus_rsp_payload_error));
  assign FetchL1Plugin_logic_banks_0_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 2'b00));
  assign FetchL1Plugin_logic_banks_0_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
  assign FetchL1Plugin_logic_banks_0_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
  assign FetchL1Plugin_logic_banks_1_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 2'b01));
  assign FetchL1Plugin_logic_banks_1_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
  assign FetchL1Plugin_logic_banks_1_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
  assign FetchL1Plugin_logic_banks_2_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 2'b10));
  assign FetchL1Plugin_logic_banks_2_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
  assign FetchL1Plugin_logic_banks_2_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
  assign FetchL1Plugin_logic_banks_3_write_valid = (FetchL1Plugin_logic_bus_rsp_valid && (FetchL1Plugin_logic_refill_onRsp_wayToAllocate == 2'b11));
  assign FetchL1Plugin_logic_banks_3_write_payload_address = {FetchL1Plugin_logic_refill_onRsp_address[11 : 6],FetchL1Plugin_logic_refill_onRsp_wordIndex};
  assign FetchL1Plugin_logic_banks_3_write_payload_data = FetchL1Plugin_logic_bus_rsp_payload_data;
  assign FetchL1Plugin_logic_bus_rsp_ready = 1'b1;
  assign when_FetchL1Plugin_l330 = (FetchL1Plugin_logic_refill_onRsp_wordIndex == 3'b111);
  assign FetchL1Plugin_logic_cmd_doIt = (fetch_logic_ctrls_1_up_ready || ((! fetch_logic_ctrls_1_up_valid) && 1'b1));
  assign FetchL1Plugin_logic_banks_0_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_0_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 3];
  assign FetchL1Plugin_logic_banks_1_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_1_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 3];
  assign FetchL1Plugin_logic_banks_2_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_2_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 3];
  assign FetchL1Plugin_logic_banks_3_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_banks_3_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 3];
  assign FetchL1Plugin_logic_ways_0_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_0_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ways_1_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_1_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ways_2_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_2_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ways_3_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_ways_3_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_plru_read_cmd_valid = FetchL1Plugin_logic_cmd_doIt;
  assign FetchL1Plugin_logic_plru_read_cmd_payload = fetch_logic_ctrls_0_down_Fetch_WORD_PC[11 : 6];
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID = (FetchL1Plugin_logic_plru_write_valid && (FetchL1Plugin_logic_plru_write_payload_address == FetchL1Plugin_logic_plru_read_cmd_payload));
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 = FetchL1Plugin_logic_plru_write_payload_data_0;
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_1 = FetchL1Plugin_logic_plru_write_payload_data_1;
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE = (|FetchL1Plugin_logic_waysWrite_mask);
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS = FetchL1Plugin_logic_waysWrite_address;
  always @(*) begin
    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_0;
    if(fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID) begin
      fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_READ_1;
    if(fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID) begin
      fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_1 = fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_1;
    end
  end

  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0 = _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1 = _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2 = _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3 = _zz_fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3;
  assign fetch_logic_ctrls_2_down_Fetch_WORD = (((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0 : 32'h0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1 : 32'h0)) | ((fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_2 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_2 : 32'h0) | (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_3 ? fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_3 : 32'h0)));
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE && (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS == fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 6]));
  assign FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_0 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[0]);
  assign FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_1 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[1]);
  assign FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_2 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[2]);
  assign FetchL1Plugin_logic_hits_w_0_indirect_translatedHits = (|{FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_2,{FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_1,FetchL1Plugin_logic_hits_w_0_indirect_wayTlbHits_0}});
  assign FetchL1Plugin_logic_hits_w_0_indirect_bypassHits = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address == _zz_FetchL1Plugin_logic_hits_w_0_indirect_bypassHits);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0 = ((fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION ? FetchL1Plugin_logic_hits_w_0_indirect_bypassHits : FetchL1Plugin_logic_hits_w_0_indirect_translatedHits) && fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded);
  assign FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_0 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[0]);
  assign FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_1 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[1]);
  assign FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_2 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[2]);
  assign FetchL1Plugin_logic_hits_w_1_indirect_translatedHits = (|{FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_2,{FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_1,FetchL1Plugin_logic_hits_w_1_indirect_wayTlbHits_0}});
  assign FetchL1Plugin_logic_hits_w_1_indirect_bypassHits = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address == _zz_FetchL1Plugin_logic_hits_w_1_indirect_bypassHits);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1 = ((fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION ? FetchL1Plugin_logic_hits_w_1_indirect_bypassHits : FetchL1Plugin_logic_hits_w_1_indirect_translatedHits) && fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded);
  assign FetchL1Plugin_logic_hits_w_2_indirect_wayTlbHits_0 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[0]);
  assign FetchL1Plugin_logic_hits_w_2_indirect_wayTlbHits_1 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[1]);
  assign FetchL1Plugin_logic_hits_w_2_indirect_wayTlbHits_2 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[2]);
  assign FetchL1Plugin_logic_hits_w_2_indirect_translatedHits = (|{FetchL1Plugin_logic_hits_w_2_indirect_wayTlbHits_2,{FetchL1Plugin_logic_hits_w_2_indirect_wayTlbHits_1,FetchL1Plugin_logic_hits_w_2_indirect_wayTlbHits_0}});
  assign FetchL1Plugin_logic_hits_w_2_indirect_bypassHits = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_address == _zz_FetchL1Plugin_logic_hits_w_2_indirect_bypassHits);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_2 = ((fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION ? FetchL1Plugin_logic_hits_w_2_indirect_bypassHits : FetchL1Plugin_logic_hits_w_2_indirect_translatedHits) && fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_loaded);
  assign FetchL1Plugin_logic_hits_w_3_indirect_wayTlbHits_0 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[0]);
  assign FetchL1Plugin_logic_hits_w_3_indirect_wayTlbHits_1 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[1]);
  assign FetchL1Plugin_logic_hits_w_3_indirect_wayTlbHits_2 = ((fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_address == fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2[31 : 12]) && fetch_logic_ctrls_1_down_MMU_WAYS_OH[2]);
  assign FetchL1Plugin_logic_hits_w_3_indirect_translatedHits = (|{FetchL1Plugin_logic_hits_w_3_indirect_wayTlbHits_2,{FetchL1Plugin_logic_hits_w_3_indirect_wayTlbHits_1,FetchL1Plugin_logic_hits_w_3_indirect_wayTlbHits_0}});
  assign FetchL1Plugin_logic_hits_w_3_indirect_bypassHits = (fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_address == _zz_FetchL1Plugin_logic_hits_w_3_indirect_bypassHits);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_3 = ((fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION ? FetchL1Plugin_logic_hits_w_3_indirect_bypassHits : FetchL1Plugin_logic_hits_w_3_indirect_translatedHits) && fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_loaded);
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT = (|{fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_3,{fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_2,{fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1,fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0}}});
  assign FetchL1Plugin_logic_ctrl_pmaPort_cmd_address = fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state = FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0[0];
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0 = (! FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_0_state);
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_1_stateSel = FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_1_state = FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_1[FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_1_stateSel];
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_1 = (! FetchL1Plugin_logic_ctrl_plruLogic_core_evict_logic_1_state);
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id = {FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_0,FetchL1Plugin_logic_ctrl_plruLogic_core_evict_sel_1};
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0[0] = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id[1];
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_update_logic_1_sel = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id[1 : 1];
  always @(*) begin
    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_1 = FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_1;
    FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_1[FetchL1Plugin_logic_ctrl_plruLogic_core_update_logic_1_sel] = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id[0];
  end

  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_0 = fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_context_state_1 = fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_1;
  assign _zz_FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id = (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 || fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_3);
  assign _zz_FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id_1 = (fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_2 || fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_3);
  assign FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id = {_zz_FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id_1,_zz_FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_id};
  always @(*) begin
    FetchL1Plugin_logic_plru_write_valid = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_valid = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_plru_write_payload_address = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_payload_address = FetchL1Plugin_logic_invalidate_counter[5:0];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_plru_write_payload_data_0 = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_payload_data_0 = _zz_FetchL1Plugin_logic_plru_write_payload_data_0[0 : 0];
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_plru_write_payload_data_1 = FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_1;
    if(when_FetchL1Plugin_l558) begin
      FetchL1Plugin_logic_plru_write_payload_data_1 = _zz_FetchL1Plugin_logic_plru_write_payload_data_0[2 : 1];
    end
  end

  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid = (fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_up_isReady);
  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address = fetch_logic_ctrls_2_down_Fetch_WORD_PC[11 : 6];
  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0 = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_0;
  assign FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_1 = FetchL1Plugin_logic_ctrl_plruLogic_core_io_update_state_1;
  assign FetchL1Plugin_logic_refill_start_wayToAllocate = FetchL1Plugin_logic_ctrl_plruLogic_core_io_evict_id;
  assign FetchL1Plugin_logic_ctrl_dataAccessFault = (_zz_FetchL1Plugin_logic_ctrl_dataAccessFault[0] && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD));
  always @(*) begin
    FetchL1Plugin_logic_trapPort_valid = 1'b0;
    if(when_FetchL1Plugin_l474) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b1;
    end
    if(when_FetchL1Plugin_l533) begin
      FetchL1Plugin_logic_trapPort_valid = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_trapPort_payload_tval = fetch_logic_ctrls_2_down_Fetch_WORD_PC;
  always @(*) begin
    FetchL1Plugin_logic_trapPort_payload_exception = 1'bx;
    if(when_FetchL1Plugin_l474) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_exception = 1'b1;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_trapPort_payload_code = 4'bxxxx;
    if(when_FetchL1Plugin_l474) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b1100;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0111;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_trapPort_payload_code = 4'b0001;
      if(when_FetchL1Plugin_l520) begin
        FetchL1Plugin_logic_trapPort_payload_code = 4'b1100;
      end
    end
  end

  assign _zz_66 = zz_FetchL1Plugin_logic_trapPort_payload_arg(1'b0);
  always @(*) FetchL1Plugin_logic_trapPort_payload_arg = _zz_66;
  always @(*) begin
    FetchL1Plugin_logic_ctrl_allowRefill = ((! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT) && (! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD));
    if(when_FetchL1Plugin_l480) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(when_FetchL1Plugin_l487) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_REFILL) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_MMU_HAZARD) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
    if(fetch_logic_ctrls_2_down_Fetch_PC_FAULT) begin
      FetchL1Plugin_logic_ctrl_allowRefill = 1'b0;
    end
  end

  assign when_FetchL1Plugin_l474 = ((! fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT) || fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD);
  assign when_FetchL1Plugin_l480 = ((FetchL1Plugin_logic_ctrl_dataAccessFault || FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault) || fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT);
  assign when_FetchL1Plugin_l487 = (fetch_logic_ctrls_2_down_MMU_PAGE_FAULT || (! fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE));
  assign when_FetchL1Plugin_l520 = (! fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION);
  always @(*) begin
    FetchL1Plugin_logic_refill_start_valid = (FetchL1Plugin_logic_ctrl_allowRefill && (! FetchL1Plugin_logic_ctrl_trapSent));
    if(when_FetchL1Plugin_l537) begin
      FetchL1Plugin_logic_refill_start_valid = 1'b0;
    end
  end

  assign FetchL1Plugin_logic_refill_start_address = fetch_logic_ctrls_2_down_MMU_TRANSLATED;
  assign FetchL1Plugin_logic_refill_start_isIo = FetchL1Plugin_logic_ctrl_pmaPort_rsp_io;
  assign fetch_logic_ctrls_2_down_TRAP = (FetchL1Plugin_logic_trapPort_valid || FetchL1Plugin_logic_ctrl_trapSent);
  assign when_FetchL1Plugin_l533 = ((! fetch_logic_ctrls_2_up_isValid) || FetchL1Plugin_logic_ctrl_trapSent);
  assign when_FetchL1Plugin_l537 = ((! fetch_logic_ctrls_2_up_isValid) && 1'b1);
  assign when_FetchL1Plugin_l541 = (((! fetch_logic_ctrls_2_up_isValid) || fetch_logic_ctrls_2_down_isReady) || fetch_logic_ctrls_2_up_isCanceling);
  assign when_FetchL1Plugin_l549 = (fetch_logic_ctrls_2_up_isValid && (! fetch_logic_ctrls_2_down_TRAP));
  assign FetchL1Plugin_logic_events_access = fetch_logic_ctrls_2_up_isMoving;
  assign FetchL1Plugin_logic_events_miss = (fetch_logic_ctrls_2_up_isMoving && FetchL1Plugin_logic_ctrl_allowRefill);
  assign FetchL1Plugin_logic_events_waiting = FetchL1Plugin_logic_ctrl_onEvents_waiting;
  assign when_FetchL1Plugin_l558 = (! FetchL1Plugin_logic_invalidate_done);
  assign _zz_FetchL1Plugin_logic_plru_write_payload_data_0 = 3'b000;
  assign LsuPlugin_logic_frontend_defaultsDecodings_0 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_1 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_2 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_3 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_4 = 1'b0;
  assign LsuPlugin_logic_frontend_defaultsDecodings_5 = 1'b0;
  always @(*) begin
    PrivilegedPlugin_logic_harts_0_xretAwayFromMachine = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        if(when_TrapPlugin_l654) begin
          PrivilegedPlugin_logic_harts_0_xretAwayFromMachine = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PrivilegedPlugin_logic_harts_0_int_pending = 1'b0;
    if(TrapPlugin_logic_harts_0_interrupt_pendingInterrupt) begin
      PrivilegedPlugin_logic_harts_0_int_pending = 1'b1;
    end
  end

  assign PrivilegedPlugin_logic_harts_0_withMachinePrivilege = (2'b11 <= PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege = (2'b01 <= PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_hartRunning = 1'b1;
  assign PrivilegedPlugin_logic_harts_0_debugMode = (! PrivilegedPlugin_logic_harts_0_hartRunning);
  always @(*) begin
    PrivilegedPlugin_logic_harts_0_m_status_sd = 1'b0;
    if(when_PrivilegedPlugin_l542) begin
      PrivilegedPlugin_logic_harts_0_m_status_sd = 1'b1;
    end
  end

  assign when_PrivilegedPlugin_l542 = (PrivilegedPlugin_logic_harts_0_m_status_fs == 2'b11);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_4 = (when_CsrService_l198 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_5 = (when_CsrService_l198 && REG_CSR_834);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_7 = (when_CsrService_l198 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_9 = (when_CsrService_l198 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_10 = (when_CsrService_l198 && REG_CSR_770);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_12 = (when_CsrService_l198 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11);
  assign _zz_when_TrapPlugin_l207 = (PrivilegedPlugin_logic_harts_0_m_ip_mtip && PrivilegedPlugin_logic_harts_0_m_ie_mtie);
  assign _zz_when_TrapPlugin_l207_1 = (PrivilegedPlugin_logic_harts_0_m_ip_msip && PrivilegedPlugin_logic_harts_0_m_ie_msie);
  assign _zz_when_TrapPlugin_l207_2 = (PrivilegedPlugin_logic_harts_0_m_ip_meip && PrivilegedPlugin_logic_harts_0_m_ie_meie);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_13 = (when_CsrService_l198 && REG_CSR_322);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_14 = (when_CsrService_l198 && _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1);
  assign PrivilegedPlugin_logic_harts_0_s_ip_seipOr = (PrivilegedPlugin_logic_harts_0_s_ip_seipSoft || PrivilegedPlugin_logic_harts_0_s_ip_seipInput);
  assign PrivilegedPlugin_logic_harts_0_s_ip_seipMasked = (PrivilegedPlugin_logic_harts_0_s_ip_seipOr && PrivilegedPlugin_logic_harts_0_m_ideleg_se);
  assign PrivilegedPlugin_logic_harts_0_s_ip_stipMasked = (PrivilegedPlugin_logic_harts_0_s_ip_stip && PrivilegedPlugin_logic_harts_0_m_ideleg_st);
  assign PrivilegedPlugin_logic_harts_0_s_ip_ssipMasked = (PrivilegedPlugin_logic_harts_0_s_ip_ssip && PrivilegedPlugin_logic_harts_0_m_ideleg_ss);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_15 = (when_CsrService_l198 && REG_CSR_260);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_16 = (when_CsrService_l198 && REG_CSR_324);
  assign _zz_when_TrapPlugin_l207_3 = (PrivilegedPlugin_logic_harts_0_s_ip_ssip && PrivilegedPlugin_logic_harts_0_s_ie_ssie);
  assign _zz_when_TrapPlugin_l207_4 = (PrivilegedPlugin_logic_harts_0_s_ip_stip && PrivilegedPlugin_logic_harts_0_s_ie_stie);
  assign _zz_when_TrapPlugin_l207_5 = (PrivilegedPlugin_logic_harts_0_s_ip_seipOr && PrivilegedPlugin_logic_harts_0_s_ie_seie);
  assign PrivilegedPlugin_logic_defaultTrap_csrPrivilege = CsrAccessPlugin_bus_decode_address[9 : 8];
  assign PrivilegedPlugin_logic_defaultTrap_csrReadOnly = (CsrAccessPlugin_bus_decode_address[11 : 10] == 2'b11);
  assign when_PrivilegedPlugin_l689 = ((PrivilegedPlugin_logic_defaultTrap_csrReadOnly && CsrAccessPlugin_bus_decode_write) || (PrivilegedPlugin_logic_harts_0_privilege < PrivilegedPlugin_logic_defaultTrap_csrPrivilege));
  assign _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH = fetch_logic_ctrls_0_down_Fetch_WORD_PC[15 : 2];
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH = ({_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[0],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[1],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[2],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[3],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[4],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH[5],{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_1,{_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_2,_zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_3}}}}}}}} ^ _zz_fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH_4);
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid = GSharePlugin_logic_mem_write_valid;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address = GSharePlugin_logic_mem_write_payload_address;
  assign fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0 = GSharePlugin_logic_mem_write_payload_data_0;
  always @(*) begin
    fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 = GSharePlugin_logic_mem_counter_spinal_port1[1 : 0];
    if(when_GSharePlugin_l88) begin
      fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0 = fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0;
    end
  end

  assign when_GSharePlugin_l88 = (fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid && (fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address == fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH));
  always @(*) begin
    BtbPlugin_logic_ras_ptr_pushIt = 1'b0;
    if(BtbPlugin_logic_applyIt_rasLogic_pushValid) begin
      BtbPlugin_logic_ras_ptr_pushIt = 1'b1;
    end
  end

  always @(*) begin
    BtbPlugin_logic_ras_ptr_popIt = 1'b0;
    if(when_BtbPlugin_l246) begin
      BtbPlugin_logic_ras_ptr_popIt = 1'b1;
    end
  end

  assign BtbPlugin_logic_ras_write_valid = BtbPlugin_logic_ras_ptr_pushIt;
  assign BtbPlugin_logic_ras_write_payload_address = BtbPlugin_logic_ras_ptr_push;
  always @(*) begin
    BtbPlugin_logic_ras_write_payload_data = 30'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    BtbPlugin_logic_ras_write_payload_data = (_zz_BtbPlugin_logic_ras_write_payload_data >>> 2'd2);
  end

  assign BtbPlugin_logic_memDp_wp_valid = BtbPlugin_logic_memWrite_valid;
  assign BtbPlugin_logic_memDp_wp_payload_address = BtbPlugin_logic_memWrite_payload_address;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_hash = BtbPlugin_logic_memWrite_payload_data_0_hash;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_pcTarget = BtbPlugin_logic_memWrite_payload_data_0_pcTarget;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_isBranch = BtbPlugin_logic_memWrite_payload_data_0_isBranch;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_isPush = BtbPlugin_logic_memWrite_payload_data_0_isPush;
  assign BtbPlugin_logic_memDp_wp_payload_data_0_isPop = BtbPlugin_logic_memWrite_payload_data_0_isPop;
  assign BtbPlugin_logic_memDp_wp_payload_mask = BtbPlugin_logic_memWrite_payload_mask;
  assign _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash = BtbPlugin_logic_mem_spinal_port1[48 : 0];
  assign BtbPlugin_logic_memDp_rp_rsp_0_hash = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[15 : 0];
  assign BtbPlugin_logic_memDp_rp_rsp_0_pcTarget = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[45 : 16];
  assign BtbPlugin_logic_memDp_rp_rsp_0_isBranch = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[46];
  assign BtbPlugin_logic_memDp_rp_rsp_0_isPush = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[47];
  assign BtbPlugin_logic_memDp_rp_rsp_0_isPop = _zz_BtbPlugin_logic_memDp_rp_rsp_0_hash[48];
  assign BtbPlugin_logic_memDp_rp_cmd_valid = BtbPlugin_logic_memRead_cmd_valid;
  assign BtbPlugin_logic_memDp_rp_cmd_payload = BtbPlugin_logic_memRead_cmd_payload;
  assign BtbPlugin_logic_memRead_rsp_0_hash = BtbPlugin_logic_memDp_rp_rsp_0_hash;
  assign BtbPlugin_logic_memRead_rsp_0_pcTarget = BtbPlugin_logic_memDp_rp_rsp_0_pcTarget;
  assign BtbPlugin_logic_memRead_rsp_0_isBranch = BtbPlugin_logic_memDp_rp_rsp_0_isBranch;
  assign BtbPlugin_logic_memRead_rsp_0_isPush = BtbPlugin_logic_memDp_rp_rsp_0_isPush;
  assign BtbPlugin_logic_memRead_rsp_0_isPop = BtbPlugin_logic_memDp_rp_rsp_0_isPop;
  assign WhiteboxerPlugin_logic_fetch_fetchId = fetch_logic_ctrls_0_down_Fetch_ID;
  assign WhiteboxerPlugin_logic_decodes_0_fire = ((decode_ctrls_0_up_LANE_SEL_0 && decode_ctrls_0_up_isReady) && (! decode_ctrls_0_lane0_upIsCancel));
  assign when_CtrlLaneApi_l50 = (decode_ctrls_0_up_isReady || decode_ctrls_0_lane0_upIsCancel);
  assign WhiteboxerPlugin_logic_decodes_0_spawn = (decode_ctrls_0_up_LANE_SEL_0 && (! decode_ctrls_0_up_LANE_SEL_0_regNext));
  assign WhiteboxerPlugin_logic_decodes_0_pc = _zz_WhiteboxerPlugin_logic_decodes_0_pc;
  assign WhiteboxerPlugin_logic_decodes_0_fetchId = decode_ctrls_0_down_Fetch_ID_0;
  assign WhiteboxerPlugin_logic_decodes_0_decodeId = decode_ctrls_0_down_Decode_DOP_ID_0;
  always @(*) begin
    early0_EnvPlugin_logic_flushPort_valid = 1'b0;
    if(when_EnvPlugin_l119) begin
      early0_EnvPlugin_logic_flushPort_valid = 1'b1;
    end
  end

  assign early0_EnvPlugin_logic_flushPort_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign early0_EnvPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    early0_EnvPlugin_logic_trapPort_valid = 1'b0;
    if(when_EnvPlugin_l119) begin
      early0_EnvPlugin_logic_trapPort_valid = 1'b1;
    end
  end

  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_exception = 1'b1;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
      end
      EnvPluginOp_ECALL : begin
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l95) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
      end
      default : begin
        if(when_EnvPlugin_l110) begin
          early0_EnvPlugin_logic_trapPort_payload_exception = 1'b0;
        end
      end
    endcase
  end

  assign early0_EnvPlugin_logic_trapPort_payload_tval = ((execute_ctrl2_down_early0_EnvPlugin_OP_lane0 == EnvPluginOp_EBREAK) ? execute_ctrl2_down_PC_lane0 : 32'h0);
  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_code = 4'b0010;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
        early0_EnvPlugin_logic_trapPort_payload_code = 4'b0011;
      end
      EnvPluginOp_ECALL : begin
        early0_EnvPlugin_logic_trapPort_payload_code = (_zz_early0_EnvPlugin_logic_trapPort_payload_code | 4'b1000);
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b0001;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l95) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b1000;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_trapPort_payload_code = 4'b0010;
      end
      default : begin
        if(when_EnvPlugin_l110) begin
          early0_EnvPlugin_logic_trapPort_payload_code = 4'b0110;
        end
      end
    endcase
  end

  always @(*) begin
    early0_EnvPlugin_logic_trapPort_payload_arg = 3'bxxx;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
      end
      EnvPluginOp_ECALL : begin
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_trapPort_payload_arg[1 : 0] = early0_EnvPlugin_logic_exe_xretPriv;
        end
      end
      EnvPluginOp_WFI : begin
      end
      EnvPluginOp_FENCE_I : begin
      end
      default : begin
      end
    endcase
  end

  assign early0_EnvPlugin_logic_exe_privilege = PrivilegedPlugin_logic_harts_0_privilege;
  assign MmuPlugin_logic_satpModeWrite = CsrAccessPlugin_bus_write_bits[31 : 31];
  assign FetchL1TileLinkPlugin_logic_down_a_valid = FetchL1Plugin_logic_bus_cmd_valid;
  assign FetchL1TileLinkPlugin_logic_down_a_payload_opcode = A_GET;
  assign FetchL1TileLinkPlugin_logic_down_a_payload_param = 3'b000;
  assign FetchL1TileLinkPlugin_logic_down_a_payload_address = FetchL1Plugin_logic_bus_cmd_payload_address;
  assign FetchL1TileLinkPlugin_logic_down_a_payload_size = 3'b110;
  assign FetchL1Plugin_logic_bus_cmd_ready = FetchL1TileLinkPlugin_logic_down_a_ready;
  assign FetchL1Plugin_logic_bus_rsp_valid = FetchL1TileLinkPlugin_logic_down_d_valid;
  assign FetchL1Plugin_logic_bus_rsp_payload_data = FetchL1TileLinkPlugin_logic_down_d_payload_data;
  assign FetchL1Plugin_logic_bus_rsp_payload_error = (FetchL1TileLinkPlugin_logic_down_d_payload_denied || FetchL1TileLinkPlugin_logic_down_d_payload_corrupt);
  assign FetchL1TileLinkPlugin_logic_down_d_ready = 1'b1;
  always @(*) begin
    DecoderPlugin_logic_forgetPort_valid = 1'b0;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_valid = 1'b1;
    end
  end

  always @(*) begin
    DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice = (decode_ctrls_1_down_PC_0 + _zz_DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice);
    end
  end

  assign PerformanceCounterPlugin_logic_commitMask = PrivilegedPlugin_logic_harts_0_commitMask;
  assign when_PerformanceCounterPlugin_l45 = (|PerformanceCounterPlugin_logic_commitMask);
  assign PerformanceCounterPlugin_logic_commitCount = (_zz_PerformanceCounterPlugin_logic_commitCount - (PerformanceCounterPlugin_logic_ignoreNextCommit && (|PerformanceCounterPlugin_logic_commitMask)));
  assign PerformanceCounterPlugin_logic_counters_cycle_needFlush = PerformanceCounterPlugin_logic_counters_cycle_value[7];
  assign PerformanceCounterPlugin_logic_counters_instret_needFlush = PerformanceCounterPlugin_logic_counters_instret_value[7];
  assign PerformanceCounterPlugin_logic_eventCycles = 1'b1;
  assign PerformanceCounterPlugin_logic_eventInstructions_0 = _zz_PerformanceCounterPlugin_logic_eventInstructions_0[0];
  always @(*) begin
    _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0)
      1'b0 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = execute_ctrl1_down_integer_RS1_lane0;
      end
      default : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = {execute_ctrl1_down_Decode_UOP_lane0[31 : 12],12'h0};
      end
    endcase
  end

  assign execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0 = _zz_execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
  always @(*) begin
    _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0)
      2'b00 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl1_down_integer_RS2_lane0;
      end
      2'b01 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = {{20{_zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0[11]}}, _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0};
      end
      2'b10 : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl1_down_PC_lane0;
      end
      default : begin
        _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = {{20{_zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1[11]}}, _zz__zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0_1};
      end
    endcase
  end

  assign execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0 = _zz_execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
  always @(*) begin
    early0_SrcPlugin_logic_addsub_combined_rs2Patched = execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0;
    if(execute_ctrl2_down_SrcStageables_REVERT_lane0) begin
      early0_SrcPlugin_logic_addsub_combined_rs2Patched = (~ execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0);
    end
    if(execute_ctrl2_down_SrcStageables_ZERO_lane0) begin
      early0_SrcPlugin_logic_addsub_combined_rs2Patched = 32'h0;
    end
  end

  assign execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0 = ($signed(_zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0) + $signed(_zz_execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0_1));
  assign execute_ctrl2_down_early0_SrcPlugin_LESS_lane0 = ((execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31] == execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[31]) ? execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0[31] : (execute_ctrl2_down_SrcStageables_UNSIGNED_lane0 ? execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0[31] : execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0[31]));
  assign lane0_IntFormatPlugin_logic_stages_0_hits = {early0_BarrelShifterPlugin_logic_wb_valid,early0_IntAluPlugin_logic_wb_valid};
  assign lane0_IntFormatPlugin_logic_stages_0_wb_valid = (execute_ctrl2_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_0_hits));
  assign lane0_IntFormatPlugin_logic_stages_0_raw = ((lane0_IntFormatPlugin_logic_stages_0_hits[0] ? early0_IntAluPlugin_logic_wb_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_0_hits[1] ? early0_BarrelShifterPlugin_logic_wb_payload : 32'h0));
  assign lane0_IntFormatPlugin_logic_stages_0_wb_payload = lane0_IntFormatPlugin_logic_stages_0_raw;
  assign lane0_IntFormatPlugin_logic_stages_1_hits = {LsuPlugin_logic_iwb_valid,early0_MulPlugin_logic_formatBus_valid};
  assign lane0_IntFormatPlugin_logic_stages_1_wb_valid = (execute_ctrl4_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_1_hits));
  assign lane0_IntFormatPlugin_logic_stages_1_raw = ((lane0_IntFormatPlugin_logic_stages_1_hits[0] ? early0_MulPlugin_logic_formatBus_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_1_hits[1] ? LsuPlugin_logic_iwb_payload : 32'h0));
  always @(*) begin
    lane0_IntFormatPlugin_logic_stages_1_wb_payload = lane0_IntFormatPlugin_logic_stages_1_raw;
    if(lane0_IntFormatPlugin_logic_stages_1_segments_0_doIt) begin
      lane0_IntFormatPlugin_logic_stages_1_wb_payload[15 : 8] = {8{lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value}};
    end
    if(lane0_IntFormatPlugin_logic_stages_1_segments_1_doIt) begin
      lane0_IntFormatPlugin_logic_stages_1_wb_payload[31 : 16] = {16{lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value}};
    end
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_1_raw[7];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value = 1'bx;
    case(execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b00 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_sels_0;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_1_segments_0_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_0_doIt = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b01);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_0 = lane0_IntFormatPlugin_logic_stages_1_raw[7];
  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_1 = lane0_IntFormatPlugin_logic_stages_1_raw[15];
  always @(*) begin
    _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = 1'bx;
    case(execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0)
      2'b00 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_0;
      end
      2'b01 : begin
        _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_sels_1;
      end
      default : begin
      end
    endcase
  end

  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 && _zz_lane0_IntFormatPlugin_logic_stages_1_segments_1_sign_value);
  assign lane0_IntFormatPlugin_logic_stages_1_segments_1_doIt = (execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 < 2'b10);
  assign lane0_IntFormatPlugin_logic_stages_2_hits = {CsrAccessPlugin_logic_wbWi_valid,early0_DivPlugin_logic_formatBus_valid};
  assign lane0_IntFormatPlugin_logic_stages_2_wb_valid = (execute_ctrl3_up_LANE_SEL_lane0 && (|lane0_IntFormatPlugin_logic_stages_2_hits));
  assign lane0_IntFormatPlugin_logic_stages_2_raw = ((lane0_IntFormatPlugin_logic_stages_2_hits[0] ? early0_DivPlugin_logic_formatBus_payload : 32'h0) | (lane0_IntFormatPlugin_logic_stages_2_hits[1] ? CsrAccessPlugin_logic_wbWi_payload : 32'h0));
  assign lane0_IntFormatPlugin_logic_stages_2_wb_payload = lane0_IntFormatPlugin_logic_stages_2_raw;
  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early0_BranchPlugin_pcCalc_target_a = execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0;
      end
      default : begin
        early0_BranchPlugin_pcCalc_target_a = execute_ctrl2_down_PC_lane0;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JAL : begin
        early0_BranchPlugin_pcCalc_target_b = {{11{_zz_early0_BranchPlugin_pcCalc_target_b[20]}}, _zz_early0_BranchPlugin_pcCalc_target_b};
      end
      BranchPlugin_BranchCtrlEnum_JALR : begin
        early0_BranchPlugin_pcCalc_target_b = {{20{_zz_early0_BranchPlugin_pcCalc_target_b_1[11]}}, _zz_early0_BranchPlugin_pcCalc_target_b_1};
      end
      default : begin
        early0_BranchPlugin_pcCalc_target_b = {{19{_zz_early0_BranchPlugin_pcCalc_target_b_2[12]}}, _zz_early0_BranchPlugin_pcCalc_target_b_2};
      end
    endcase
  end

  assign early0_BranchPlugin_pcCalc_slices = (_zz_early0_BranchPlugin_pcCalc_slices + {1'b0,1'b1});
  always @(*) begin
    execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
    execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[0] = 1'b0;
  end

  assign execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = (execute_ctrl2_down_PC_lane0 + _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = (execute_ctrl2_down_PC_lane0 + _zz_execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0);
  assign AlignerPlugin_logic_maskGen_frontMasks_0 = 1'b1;
  assign AlignerPlugin_logic_maskGen_backMasks_0 = 1'b1;
  assign fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK = (AlignerPlugin_logic_maskGen_frontMasks_0 & ((! fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED) ? 1'b1 : AlignerPlugin_logic_maskGen_backMasks_0));
  assign fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_LAST = ((fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED) ? 1'b1 : 1'b0);
  assign AlignerPlugin_logic_slicesInstructions_0 = AlignerPlugin_logic_slices_data_0;
  always @(*) begin
    AlignerPlugin_logic_scanners_0_usageMask = 1'b0;
    AlignerPlugin_logic_scanners_0_usageMask[0] = AlignerPlugin_logic_scanners_0_checker_0_required;
  end

  assign AlignerPlugin_logic_scanners_0_checker_0_required = 1'b1;
  assign AlignerPlugin_logic_scanners_0_checker_0_last = (AlignerPlugin_logic_slices_data_0[1 : 0] != 2'b11);
  assign AlignerPlugin_logic_scanners_0_checker_0_redo = 1'b0;
  assign AlignerPlugin_logic_scanners_0_checker_0_present = AlignerPlugin_logic_slices_mask[0];
  assign AlignerPlugin_logic_scanners_0_checker_0_valid = AlignerPlugin_logic_scanners_0_checker_0_present;
  assign AlignerPlugin_logic_scanners_0_redo = (|AlignerPlugin_logic_scanners_0_checker_0_redo);
  assign AlignerPlugin_logic_scanners_0_valid = (AlignerPlugin_logic_scanners_0_checker_0_valid && (1'b1 || (|AlignerPlugin_logic_scanners_0_checker_0_redo)));
  assign AlignerPlugin_logic_usedMask_0 = 1'b0;
  assign AlignerPlugin_logic_extractors_0_first = 1'b1;
  assign AlignerPlugin_logic_extractors_0_usableMask = (AlignerPlugin_logic_scanners_0_valid && (! AlignerPlugin_logic_usedMask_0[0]));
  assign AlignerPlugin_logic_extractors_0_usableMask_bools_0 = AlignerPlugin_logic_extractors_0_usableMask[0];
  assign _zz_AlignerPlugin_logic_extractors_0_slicesOh[0] = (AlignerPlugin_logic_extractors_0_usableMask_bools_0 && (! 1'b0));
  assign AlignerPlugin_logic_extractors_0_slicesOh = _zz_AlignerPlugin_logic_extractors_0_slicesOh;
  always @(*) begin
    AlignerPlugin_logic_extractors_0_redo = AlignerPlugin_logic_scanners_0_redo;
    if(when_AlignerPlugin_l160) begin
      AlignerPlugin_logic_extractors_0_redo = 1'b0;
    end
  end

  assign AlignerPlugin_logic_extractors_0_localMask = AlignerPlugin_logic_scanners_0_checker_0_required;
  always @(*) begin
    AlignerPlugin_logic_extractors_0_usageMask = AlignerPlugin_logic_scanners_0_usageMask;
    if(when_AlignerPlugin_l160) begin
      AlignerPlugin_logic_extractors_0_usageMask = 1'b0;
    end
  end

  assign AlignerPlugin_logic_usedMask_1 = (AlignerPlugin_logic_usedMask_0 | AlignerPlugin_logic_extractors_0_usageMask);
  always @(*) begin
    AlignerPlugin_logic_extractors_0_valid = (|AlignerPlugin_logic_extractors_0_slicesOh);
    if(when_AlignerPlugin_l160) begin
      AlignerPlugin_logic_extractors_0_valid = 1'b0;
    end
  end

  assign when_AlignerPlugin_l160 = (AlignerPlugin_api_haltIt || (AlignerPlugin_api_singleFetch && (! AlignerPlugin_logic_extractors_0_first)));
  assign when_AlignerPlugin_l171 = (decode_ctrls_0_up_isFiring && 1'b1);
  assign AlignerPlugin_logic_feeder_lanes_0_valid = AlignerPlugin_logic_extractors_0_valid;
  assign decode_ctrls_0_up_LANE_SEL_0 = AlignerPlugin_logic_feeder_lanes_0_valid;
  assign decode_ctrls_0_up_Decode_INSTRUCTION_0 = AlignerPlugin_logic_extractors_0_ctx_instruction;
  assign decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0 = 1'b0;
  always @(*) begin
    decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0 = AlignerPlugin_logic_extractors_0_ctx_instruction;
    if(AlignerPlugin_logic_feeder_lanes_0_isRvc) begin
      decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0[31 : 16] = 16'h0;
    end
  end

  assign AlignerPlugin_logic_feeder_lanes_0_isRvc = (AlignerPlugin_logic_extractors_0_ctx_instruction[1 : 0] != 2'b11);
  assign decode_ctrls_0_up_PC_0 = AlignerPlugin_logic_extractors_0_ctx_pc;
  assign decode_ctrls_0_up_Decode_DOP_ID_0 = AlignerPlugin_logic_feeder_harts_0_dopId;
  assign decode_ctrls_0_up_Fetch_ID_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID;
  assign decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0 = AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY;
  assign decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH;
  assign decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN;
  assign decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC;
  assign decode_ctrls_0_up_Prediction_WORD_JUMPED_0 = AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED;
  assign decode_ctrls_0_up_TRAP_0 = AlignerPlugin_logic_extractors_0_ctx_trap;
  assign AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction = 1'b1;
  assign decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0 = (decode_ctrls_0_up_Prediction_WORD_JUMPED_0 && AlignerPlugin_logic_feeder_lanes_0_onBtb_didPrediction);
  assign decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0 = decode_ctrls_0_up_Prediction_WORD_JUMP_PC_0;
  assign decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0 = decode_ctrls_0_up_Prediction_WORD_SLICES_BRANCH_0;
  assign decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0 = decode_ctrls_0_up_Prediction_WORD_SLICES_TAKEN_0;
  assign decode_ctrls_0_up_Prediction_ALIGN_REDO_0 = AlignerPlugin_logic_extractors_0_redo;
  assign decode_ctrls_0_up_valid = (|AlignerPlugin_logic_feeder_lanes_0_valid);
  assign AlignerPlugin_logic_nobuffer_remaningMask = (AlignerPlugin_logic_nobuffer_mask & (~ AlignerPlugin_logic_usedMask_1));
  assign when_AlignerPlugin_l292 = (decode_ctrls_0_up_isValid && decode_ctrls_0_up_isReady);
  assign CfuPlugin_logic_onFork_functionsIds_0 = execute_ctrl2_down_Decode_UOP_lane0[14 : 12];
  assign CfuPlugin_logic_onFork_functionsIds_1 = execute_ctrl2_down_Decode_UOP_lane0[14 : 12];
  assign CfuPlugin_logic_bus_cmd_payload_cfu_index = CfuPlugin_logic_csr_cfuIndex;
  assign CfuPlugin_logic_bus_cmd_payload_state_index = CfuPlugin_logic_csr_stateId;
  assign CfuPlugin_logic_bus_cmd_payload_function_id = _zz_CfuPlugin_logic_bus_cmd_payload_function_id;
  assign CfuPlugin_logic_bus_cmd_payload_raw_insn = execute_ctrl2_down_Decode_UOP_lane0;
  assign CfuPlugin_logic_bus_cmd_payload_inputs_0 = execute_ctrl2_up_integer_RS1_lane0;
  always @(*) begin
    case(execute_ctrl2_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0)
      Input2Kind_RS : begin
        _zz_CfuPlugin_logic_bus_cmd_payload_inputs_1 = execute_ctrl2_up_integer_RS2_lane0;
      end
      default : begin
        _zz_CfuPlugin_logic_bus_cmd_payload_inputs_1 = _zz__zz_CfuPlugin_logic_bus_cmd_payload_inputs_1;
      end
    endcase
  end

  assign CfuPlugin_logic_bus_cmd_payload_inputs_1 = _zz_CfuPlugin_logic_bus_cmd_payload_inputs_1;
  assign CfuPlugin_logic_bus_rsp_ready = 1'b1;
  assign CfuPlugin_logic_bus_rsp_toFlow_valid = CfuPlugin_logic_bus_rsp_valid;
  assign CfuPlugin_logic_bus_rsp_toFlow_payload_outputs_0 = CfuPlugin_logic_bus_rsp_payload_outputs_0;
  assign CfuPlugin_logic_onJoin_busRspStream_valid = CfuPlugin_logic_bus_rsp_toFlow_valid;
  assign CfuPlugin_logic_onJoin_busRspStream_payload_outputs_0 = CfuPlugin_logic_bus_rsp_toFlow_payload_outputs_0;
  assign CfuPlugin_logic_onJoin_busRspStream_ready = CfuPlugin_logic_onJoin_busRspStream_fifo_io_push_ready;
  assign CfuPlugin_logic_onJoin_freezeIt = (execute_ctrl4_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0 && (! CfuPlugin_logic_onJoin_busRspStream_fifo_io_pop_valid));
  assign CfuPlugin_logic_onJoin_busRspStream_fifo_io_pop_ready = (execute_ctrl4_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0 && (! execute_freeze_valid));
  assign CfuPlugin_logic_wb_valid = (execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_CfuPlugin_logic_CFU_ENABLE_lane0);
  assign CfuPlugin_logic_wb_payload = CfuPlugin_logic_onJoin_busRspStream_fifo_io_pop_payload_outputs_0;
  assign execute_ctrl0_down_AguPlugin_SIZE_lane0 = execute_ctrl0_down_Decode_UOP_lane0[13 : 12];
  assign LsuPlugin_logic_flusher_wantExit = 1'b0;
  always @(*) begin
    LsuPlugin_logic_flusher_wantStart = 1'b0;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_CMD : begin
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
      end
      default : begin
        LsuPlugin_logic_flusher_wantStart = 1'b1;
      end
    endcase
  end

  assign LsuPlugin_logic_flusher_wantKill = 1'b0;
  assign TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready = LsuPlugin_logic_flusher_arbiter_io_inputs_0_ready;
  assign LsuPlugin_logic_flusher_inflight = (|{(execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuL1_FLUSH_lane0),(execute_ctrl3_down_LsuL1_SEL_lane0 && execute_ctrl3_down_LsuL1_FLUSH_lane0)});
  assign early0_EnvPlugin_logic_exe_xretPriv = execute_ctrl2_down_Decode_UOP_lane0[29 : 28];
  always @(*) begin
    early0_EnvPlugin_logic_exe_commit = 1'b0;
    case(execute_ctrl2_down_early0_EnvPlugin_OP_lane0)
      EnvPluginOp_EBREAK : begin
      end
      EnvPluginOp_ECALL : begin
      end
      EnvPluginOp_PRIV_RET : begin
        if(when_EnvPlugin_l86) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
      EnvPluginOp_WFI : begin
        if(when_EnvPlugin_l95) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
      EnvPluginOp_FENCE_I : begin
        early0_EnvPlugin_logic_exe_commit = 1'b1;
      end
      default : begin
        if(when_EnvPlugin_l110) begin
          early0_EnvPlugin_logic_exe_commit = 1'b1;
        end
      end
    endcase
  end

  assign early0_EnvPlugin_logic_exe_retKo = ((PrivilegedPlugin_logic_harts_0_m_status_tsr && (early0_EnvPlugin_logic_exe_privilege == 2'b01)) && (early0_EnvPlugin_logic_exe_xretPriv == 2'b01));
  assign early0_EnvPlugin_logic_exe_vmaKo = (((early0_EnvPlugin_logic_exe_privilege == 2'b01) && PrivilegedPlugin_logic_harts_0_m_status_tvm) || (early0_EnvPlugin_logic_exe_privilege == 2'b00));
  assign when_EnvPlugin_l86 = ((early0_EnvPlugin_logic_exe_xretPriv <= PrivilegedPlugin_logic_harts_0_privilege) && (! early0_EnvPlugin_logic_exe_retKo));
  assign when_EnvPlugin_l95 = ((early0_EnvPlugin_logic_exe_privilege == 2'b11) || ((! PrivilegedPlugin_logic_harts_0_m_status_tw) && (1'b0 || (early0_EnvPlugin_logic_exe_privilege == 2'b01))));
  assign when_EnvPlugin_l110 = (! early0_EnvPlugin_logic_exe_vmaKo);
  assign when_EnvPlugin_l119 = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_early0_EnvPlugin_SEL_lane0);
  assign when_EnvPlugin_l123 = (! early0_EnvPlugin_logic_exe_commit);
  assign execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0 = ($signed(execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0) == $signed(execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0));
  assign execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 = (execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0 != execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0);
  assign early0_BranchPlugin_logic_alu_expectedMsb = (MmuPlugin_api_fetchTranslationEnable ? _zz_early0_BranchPlugin_logic_alu_expectedMsb[31] : 1'b0);
  assign execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = ((execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR) && 1'b0);
  assign switch_Misc_l242 = execute_ctrl3_down_Decode_UOP_lane0[14 : 12];
  always @(*) begin
    casez(switch_Misc_l242)
      3'b000 : begin
        _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = execute_ctrl3_down_early0_BranchPlugin_logic_alu_EQ_lane0;
      end
      3'b001 : begin
        _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! execute_ctrl3_down_early0_BranchPlugin_logic_alu_EQ_lane0);
      end
      3'b1?1 : begin
        _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = (! execute_ctrl3_down_early0_SrcPlugin_LESS_lane0);
      end
      default : begin
        _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = execute_ctrl3_down_early0_SrcPlugin_LESS_lane0;
      end
    endcase
  end

  always @(*) begin
    case(execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0)
      BranchPlugin_BranchCtrlEnum_JALR : begin
        _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      BranchPlugin_BranchCtrlEnum_JAL : begin
        _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = 1'b1;
      end
      default : begin
        _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1 = _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
      end
    endcase
  end

  assign execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 = _zz_execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0_1;
  assign execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0 = (execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 ? execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 : execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_wrongCond = (execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0 != execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_needFix = ((early0_BranchPlugin_logic_jumpLogic_wrongCond || (execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0 && execute_ctrl3_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0)) || execute_ctrl3_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0);
  assign early0_BranchPlugin_logic_jumpLogic_doIt = ((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_down_early0_BranchPlugin_SEL_lane0) && early0_BranchPlugin_logic_jumpLogic_needFix);
  assign early0_BranchPlugin_logic_jumpLogic_history_shifter = execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
  assign when_BranchPlugin_l218 = (execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign early0_BranchPlugin_logic_jumpLogic_history_next = early0_BranchPlugin_logic_jumpLogic_history_shifter_1;
  assign early0_BranchPlugin_logic_jumpLogic_history_fetched = execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
  assign early0_BranchPlugin_logic_pcPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_pcPort_payload_fault = execute_ctrl3_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  assign early0_BranchPlugin_logic_pcPort_payload_pc = execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_btb_REAL_TARGET_lane0;
  assign early0_BranchPlugin_logic_historyPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_historyPort_payload_history = early0_BranchPlugin_logic_jumpLogic_history_next;
  assign early0_BranchPlugin_logic_flushPort_valid = early0_BranchPlugin_logic_jumpLogic_doIt;
  assign early0_BranchPlugin_logic_flushPort_payload_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign early0_BranchPlugin_logic_flushPort_payload_self = 1'b0;
  assign execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0 = ((execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0[1 : 0] != 2'b00) && execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0);
  always @(*) begin
    early0_BranchPlugin_logic_trapPort_valid = 1'b0;
    if(when_BranchPlugin_l251) begin
      early0_BranchPlugin_logic_trapPort_valid = 1'b1;
    end
  end

  assign early0_BranchPlugin_logic_trapPort_payload_exception = 1'b1;
  assign early0_BranchPlugin_logic_trapPort_payload_code = 4'b0000;
  assign early0_BranchPlugin_logic_trapPort_payload_tval = execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign early0_BranchPlugin_logic_trapPort_payload_arg = 3'b000;
  assign when_BranchPlugin_l251 = (early0_BranchPlugin_logic_jumpLogic_doIt && execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_MISSALIGNED_lane0);
  assign execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 = (execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JAL);
  assign execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 = (execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_JALR);
  assign early0_BranchPlugin_logic_jumpLogic_rdLink = (|{(execute_ctrl3_down_Decode_UOP_lane0[11 : 7] == 5'h05),(execute_ctrl3_down_Decode_UOP_lane0[11 : 7] == 5'h01)});
  assign early0_BranchPlugin_logic_jumpLogic_rs1Link = (|{(execute_ctrl3_down_Decode_UOP_lane0[19 : 15] == 5'h05),(execute_ctrl3_down_Decode_UOP_lane0[19 : 15] == 5'h01)});
  assign early0_BranchPlugin_logic_jumpLogic_rdEquRs1 = (execute_ctrl3_down_Decode_UOP_lane0[11 : 7] == execute_ctrl3_down_Decode_UOP_lane0[19 : 15]);
  assign early0_BranchPlugin_logic_jumpLogic_learn_valid = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_down_isReady) && (! execute_lane0_ctrls_3_upIsCancel)) && (|execute_ctrl3_down_early0_BranchPlugin_SEL_lane0));
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_taken = execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_COND_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget = execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice = execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch = (execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 == BranchPlugin_BranchCtrlEnum_B);
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_isPush = ((execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JAL_lane0 || execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0) && early0_BranchPlugin_logic_jumpLogic_rdLink);
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_isPop = (execute_ctrl3_down_early0_BranchPlugin_logic_jumpLogic_IS_JALR_lane0 && (((! early0_BranchPlugin_logic_jumpLogic_rdLink) && early0_BranchPlugin_logic_jumpLogic_rs1Link) || ((early0_BranchPlugin_logic_jumpLogic_rdLink && early0_BranchPlugin_logic_jumpLogic_rs1Link) && (! early0_BranchPlugin_logic_jumpLogic_rdEquRs1))));
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong = early0_BranchPlugin_logic_jumpLogic_needFix;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget = execute_ctrl3_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_history = early0_BranchPlugin_logic_jumpLogic_history_fetched;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign early0_BranchPlugin_logic_events_branchMiss = ((early0_BranchPlugin_logic_jumpLogic_learn_valid && early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch) && early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong);
  assign early0_BranchPlugin_logic_events_branchCount = (early0_BranchPlugin_logic_jumpLogic_learn_valid && early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch);
  assign early0_BranchPlugin_logic_wb_valid = execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
  assign early0_BranchPlugin_logic_wb_payload = execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign execute_ctrl2_COMPLETED_lane0_bypass = (execute_ctrl2_up_COMPLETED_lane0 || execute_ctrl2_down_COMPLETION_AT_2_lane0);
  assign execute_ctrl3_COMPLETED_lane0_bypass = (execute_ctrl3_up_COMPLETED_lane0 || execute_ctrl3_down_COMPLETION_AT_3_lane0);
  assign execute_ctrl4_COMPLETED_lane0_bypass = (execute_ctrl4_up_COMPLETED_lane0 || execute_ctrl4_down_COMPLETION_AT_4_lane0);
  assign execute_lane0_api_hartsInflight[0] = (|{(execute_ctrl4_up_LANE_SEL_lane0 && 1'b1),{(execute_ctrl3_up_LANE_SEL_lane0 && 1'b1),{(execute_ctrl2_up_LANE_SEL_lane0 && 1'b1),(execute_ctrl1_up_LANE_SEL_lane0 && 1'b1)}}});
  assign LearnPlugin_logic_buffered_0_valid = early0_BranchPlugin_logic_jumpLogic_learn_valid;
  assign early0_BranchPlugin_logic_jumpLogic_learn_ready = LearnPlugin_logic_buffered_0_ready;
  assign LearnPlugin_logic_buffered_0_payload_pcOnLastSlice = early0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  assign LearnPlugin_logic_buffered_0_payload_pcTarget = early0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  assign LearnPlugin_logic_buffered_0_payload_taken = early0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  assign LearnPlugin_logic_buffered_0_payload_isBranch = early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  assign LearnPlugin_logic_buffered_0_payload_isPush = early0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  assign LearnPlugin_logic_buffered_0_payload_isPop = early0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  assign LearnPlugin_logic_buffered_0_payload_wasWrong = early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  assign LearnPlugin_logic_buffered_0_payload_badPredictedTarget = early0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  assign LearnPlugin_logic_buffered_0_payload_history = early0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  assign LearnPlugin_logic_buffered_0_payload_uopId = early0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  assign LearnPlugin_logic_buffered_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_buffered_0_ready = streamArbiter_10_io_inputs_0_ready;
  assign LearnPlugin_logic_arbitrated_valid = streamArbiter_10_io_output_valid;
  assign LearnPlugin_logic_arbitrated_payload_pcOnLastSlice = streamArbiter_10_io_output_payload_pcOnLastSlice;
  assign LearnPlugin_logic_arbitrated_payload_pcTarget = streamArbiter_10_io_output_payload_pcTarget;
  assign LearnPlugin_logic_arbitrated_payload_taken = streamArbiter_10_io_output_payload_taken;
  assign LearnPlugin_logic_arbitrated_payload_isBranch = streamArbiter_10_io_output_payload_isBranch;
  assign LearnPlugin_logic_arbitrated_payload_isPush = streamArbiter_10_io_output_payload_isPush;
  assign LearnPlugin_logic_arbitrated_payload_isPop = streamArbiter_10_io_output_payload_isPop;
  assign LearnPlugin_logic_arbitrated_payload_wasWrong = streamArbiter_10_io_output_payload_wasWrong;
  assign LearnPlugin_logic_arbitrated_payload_badPredictedTarget = streamArbiter_10_io_output_payload_badPredictedTarget;
  assign LearnPlugin_logic_arbitrated_payload_history = streamArbiter_10_io_output_payload_history;
  assign LearnPlugin_logic_arbitrated_payload_uopId = streamArbiter_10_io_output_payload_uopId;
  assign LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = streamArbiter_10_io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_arbitrated_ready = 1'b1;
  assign LearnPlugin_logic_arbitrated_toFlow_valid = LearnPlugin_logic_arbitrated_valid;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_pcOnLastSlice = LearnPlugin_logic_arbitrated_payload_pcOnLastSlice;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_pcTarget = LearnPlugin_logic_arbitrated_payload_pcTarget;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_taken = LearnPlugin_logic_arbitrated_payload_taken;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_isBranch = LearnPlugin_logic_arbitrated_payload_isBranch;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_isPush = LearnPlugin_logic_arbitrated_payload_isPush;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_isPop = LearnPlugin_logic_arbitrated_payload_isPop;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_wasWrong = LearnPlugin_logic_arbitrated_payload_wasWrong;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_badPredictedTarget = LearnPlugin_logic_arbitrated_payload_badPredictedTarget;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_history = LearnPlugin_logic_arbitrated_payload_history;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_uopId = LearnPlugin_logic_arbitrated_payload_uopId;
  assign LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = LearnPlugin_logic_arbitrated_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign LearnPlugin_logic_learn_valid = LearnPlugin_logic_arbitrated_toFlow_valid;
  assign LearnPlugin_logic_learn_payload_pcOnLastSlice = LearnPlugin_logic_arbitrated_toFlow_payload_pcOnLastSlice;
  assign LearnPlugin_logic_learn_payload_pcTarget = LearnPlugin_logic_arbitrated_toFlow_payload_pcTarget;
  assign LearnPlugin_logic_learn_payload_taken = LearnPlugin_logic_arbitrated_toFlow_payload_taken;
  assign LearnPlugin_logic_learn_payload_isBranch = LearnPlugin_logic_arbitrated_toFlow_payload_isBranch;
  assign LearnPlugin_logic_learn_payload_isPush = LearnPlugin_logic_arbitrated_toFlow_payload_isPush;
  assign LearnPlugin_logic_learn_payload_isPop = LearnPlugin_logic_arbitrated_toFlow_payload_isPop;
  assign LearnPlugin_logic_learn_payload_wasWrong = LearnPlugin_logic_arbitrated_toFlow_payload_wasWrong;
  assign LearnPlugin_logic_learn_payload_badPredictedTarget = LearnPlugin_logic_arbitrated_toFlow_payload_badPredictedTarget;
  assign LearnPlugin_logic_learn_payload_history = LearnPlugin_logic_arbitrated_toFlow_payload_history;
  assign LearnPlugin_logic_learn_payload_uopId = LearnPlugin_logic_arbitrated_toFlow_payload_uopId;
  assign LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = LearnPlugin_logic_arbitrated_toFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign when_DecoderPlugin_l143 = (decode_ctrls_1_up_isMoving && 1'b1);
  assign DecoderPlugin_logic_interrupt_async = PrivilegedPlugin_logic_harts_0_int_pending;
  assign when_DecoderPlugin_l151 = (((! decode_ctrls_1_up_valid) || decode_ctrls_1_up_ready) || decode_ctrls_1_up_isCanceling);
  assign _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00000018) == 32'h0);
  assign decode_ctrls_1_down_RS1_ENABLE_0 = _zz_decode_ctrls_1_down_RS1_ENABLE_0[0];
  assign decode_ctrls_1_down_RS1_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[19 : 15];
  assign decode_ctrls_1_down_RS2_ENABLE_0 = _zz_decode_ctrls_1_down_RS2_ENABLE_0[0];
  assign decode_ctrls_1_down_RS2_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[24 : 20];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000000c) == 32'h00000008);
  always @(*) begin
    decode_ctrls_1_down_RD_ENABLE_0 = _zz_decode_ctrls_1_down_RD_ENABLE_0[0];
    if(when_DecoderPlugin_l247) begin
      decode_ctrls_1_down_RD_ENABLE_0 = 1'b0;
    end
  end

  assign decode_ctrls_1_down_RD_PHYS_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0[11 : 7];
  always @(*) begin
    decode_ctrls_1_down_Decode_LEGAL_0 = ((|{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000005f) == 32'h00000017),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0000005f) == 32'h0000000b),{((decode_ctrls_1_down_Decode_INSTRUCTION_0 & _zz_decode_ctrls_1_down_Decode_LEGAL_0) == 32'h0000006f),{(_zz_decode_ctrls_1_down_Decode_LEGAL_0_1 == _zz_decode_ctrls_1_down_Decode_LEGAL_0_2),{_zz_decode_ctrls_1_down_Decode_LEGAL_0_3,{_zz_decode_ctrls_1_down_Decode_LEGAL_0_4,_zz_decode_ctrls_1_down_Decode_LEGAL_0_5}}}}}}) && (! decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0));
    if(when_CfuPlugin_l115) begin
      decode_ctrls_1_down_Decode_LEGAL_0 = 1'b0;
    end
  end

  assign when_CfuPlugin_l115 = (decode_ctrls_1_down_CfuPlugin_logic_CFU_ENABLE_0 && (! CfuPlugin_logic_en));
  assign DecoderPlugin_logic_laneLogic_0_interruptPending = DecoderPlugin_logic_interrupt_buffered[0];
  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_valid = 1'b0;
    if(when_DecoderPlugin_l229) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_valid = ((! decode_ctrls_1_up_TRAP_0) || DecoderPlugin_logic_laneLogic_0_interruptPending);
      if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
        DecoderPlugin_logic_laneLogic_0_trapPort_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b1;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b0;
    end
    if(DecoderPlugin_logic_laneLogic_0_interruptPending) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception = 1'b0;
    end
  end

  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval = decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0;
  always @(*) begin
    DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0010;
    if(DecoderPlugin_logic_laneLogic_0_fixer_doIt) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0100;
    end
    if(DecoderPlugin_logic_laneLogic_0_interruptPending) begin
      DecoderPlugin_logic_laneLogic_0_trapPort_payload_code = 4'b0000;
    end
  end

  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_laneAge = 1'b0;
  assign DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg = 3'b000;
  assign DecoderPlugin_logic_laneLogic_0_fixer_isJb = _zz_DecoderPlugin_logic_laneLogic_0_fixer_isJb[0];
  assign DecoderPlugin_logic_laneLogic_0_fixer_doIt = (decode_ctrls_1_up_LANE_SEL_0 && ((decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0 && (! DecoderPlugin_logic_laneLogic_0_fixer_isJb)) || decode_ctrls_1_down_Prediction_ALIGN_REDO_0));
  assign when_CtrlLaneApi_l50_1 = (decode_ctrls_1_up_isReady || decode_ctrls_1_lane0_upIsCancel);
  assign DecoderPlugin_logic_laneLogic_0_completionPort_valid = ((decode_ctrls_1_up_LANE_SEL_0 && decode_ctrls_1_down_TRAP_0) && (decode_ctrls_1_up_LANE_SEL_0 && (! decode_ctrls_1_up_LANE_SEL_0_regNext)));
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap = 1'b1;
  assign DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit = 1'b0;
  assign when_DecoderPlugin_l229 = (decode_ctrls_1_up_LANE_SEL_0 && (((! decode_ctrls_1_down_Decode_LEGAL_0) || DecoderPlugin_logic_laneLogic_0_interruptPending) || DecoderPlugin_logic_laneLogic_0_fixer_doIt));
  assign DecoderPlugin_logic_laneLogic_0_flushPort_valid = (decode_ctrls_1_up_LANE_SEL_0 && decode_ctrls_1_down_TRAP_0);
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DecoderPlugin_logic_laneLogic_0_flushPort_payload_self = 1'b0;
  assign when_DecoderPlugin_l247 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0[11 : 7] == 5'h0) && (|1'b1));
  assign decode_ctrls_1_down_Decode_UOP_0 = decode_ctrls_1_down_Decode_INSTRUCTION_0;
  assign DecoderPlugin_logic_laneLogic_0_uopIdBase = DecoderPlugin_logic_harts_0_uopId;
  assign decode_ctrls_1_down_Decode_UOP_ID_0 = (DecoderPlugin_logic_laneLogic_0_uopIdBase + 16'h0);
  assign DispatchPlugin_logic_trapPendings[0] = 1'b0;
  assign DispatchPlugin_logic_candidates_0_moving = (((! DispatchPlugin_logic_candidates_0_ctx_valid) || DispatchPlugin_logic_candidates_0_fire) || DispatchPlugin_logic_candidates_0_cancel);
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && 1'b1) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS)) && 1'b1) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))}));
  assign DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard = (DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE && (|{((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && 1'b1) && (! execute_ctrl2_down_BYPASSED_AT_3_lane0)),((((DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 && execute_ctrl1_up_RD_ENABLE_lane0) && (execute_ctrl1_up_RD_PHYS_lane0 == DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS)) && 1'b1) && (! execute_ctrl1_down_BYPASSED_AT_2_lane0))}));
  assign DispatchPlugin_logic_candidates_0_rsHazards[0] = (|{DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_1_hazard,DispatchPlugin_logic_rsHazardChecker_0_onLl_0_onRs_0_hazard});
  assign DispatchPlugin_logic_reservationChecker_0_onLl_0_hit = 1'b0;
  assign DispatchPlugin_logic_candidates_0_reservationHazards[0] = DispatchPlugin_logic_reservationChecker_0_onLl_0_hit;
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0 = (|{(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0),(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl1_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0)});
  assign DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1 = (|(((DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 && execute_ctrl2_up_LANE_SEL_lane0) && 1'b1) && execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0));
  assign DispatchPlugin_logic_flushChecker_0_oldersHazard = 1'b0;
  assign DispatchPlugin_logic_candidates_0_flushHazards = ((|{DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_1,DispatchPlugin_logic_flushChecker_0_executeCheck_0_hits_0}) || (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES && DispatchPlugin_logic_flushChecker_0_oldersHazard));
  assign DispatchPlugin_logic_fenceChecker_olderInflights = (|execute_lane0_api_hartsInflight[0]);
  assign DispatchPlugin_logic_candidates_0_fenceOlderHazards = (DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER && (DispatchPlugin_logic_fenceChecker_olderInflights[0] || 1'b0));
  always @(*) begin
    decode_ctrls_1_down_ready = 1'b1;
    if(when_DispatchPlugin_l368) begin
      decode_ctrls_1_down_ready = 1'b0;
    end
  end

  assign DispatchPlugin_logic_feeds_0_sending = DispatchPlugin_logic_candidates_0_fire;
  assign DispatchPlugin_logic_candidates_0_cancel = decode_ctrls_1_lane0_upIsCancel;
  assign DispatchPlugin_logic_candidates_0_ctx_valid = ((decode_ctrls_1_up_isValid && decode_ctrls_1_up_LANE_SEL_0) && (! DispatchPlugin_logic_feeds_0_sent));
  always @(*) begin
    DispatchPlugin_logic_candidates_0_ctx_laneLayerHits = decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0;
    if(decode_ctrls_1_down_TRAP_0) begin
      DispatchPlugin_logic_candidates_0_ctx_laneLayerHits = 1'b1;
    end
  end

  assign DispatchPlugin_logic_candidates_0_ctx_uop = decode_ctrls_1_down_Decode_UOP_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED = decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC = decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN = decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH = decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY = decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER = decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH = decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH = decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES = decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3 = decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4 = decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_PC = decode_ctrls_1_down_PC_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_TRAP = decode_ctrls_1_down_TRAP_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE = decode_ctrls_1_down_RS1_ENABLE_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS = decode_ctrls_1_down_RS1_PHYS_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE = decode_ctrls_1_down_RS2_ENABLE_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS = decode_ctrls_1_down_RS2_PHYS_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE = decode_ctrls_1_down_RD_ENABLE_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS = decode_ctrls_1_down_RD_PHYS_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0;
  assign DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0 = decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0;
  assign when_DispatchPlugin_l368 = ((decode_ctrls_1_up_LANE_SEL_0 && (! DispatchPlugin_logic_feeds_0_sent)) && (! DispatchPlugin_logic_candidates_0_fire));
  assign DispatchPlugin_logic_scheduler_eusFree_0 = 1'b1;
  assign DispatchPlugin_logic_scheduler_hartFree_0 = 1'b1;
  assign DispatchPlugin_logic_scheduler_arbiters_0_candHazard = 1'b0;
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits = (((DispatchPlugin_logic_candidates_0_ctx_laneLayerHits & (~ DispatchPlugin_logic_candidates_0_rsHazards)) & (~ DispatchPlugin_logic_candidates_0_reservationHazards)) & DispatchPlugin_logic_scheduler_eusFree_0[0]);
  assign DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 = DispatchPlugin_logic_scheduler_arbiters_0_layersHits[0];
  assign _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh[0] = (DispatchPlugin_logic_scheduler_arbiters_0_layersHits_bools_0 && (! 1'b0));
  assign DispatchPlugin_logic_scheduler_arbiters_0_layerOh = _zz_DispatchPlugin_logic_scheduler_arbiters_0_layerOh;
  assign DispatchPlugin_logic_scheduler_arbiters_0_eusOh = (|DispatchPlugin_logic_scheduler_arbiters_0_layerOh[0]);
  assign DispatchPlugin_logic_scheduler_arbiters_0_doIt = (((((DispatchPlugin_logic_candidates_0_ctx_valid && (! DispatchPlugin_logic_candidates_0_flushHazards)) && (! DispatchPlugin_logic_candidates_0_fenceOlderHazards)) && (|DispatchPlugin_logic_scheduler_arbiters_0_layerOh)) && DispatchPlugin_logic_scheduler_hartFree_0[0]) && (! DispatchPlugin_logic_scheduler_arbiters_0_candHazard));
  assign DispatchPlugin_logic_scheduler_eusFree_1 = (DispatchPlugin_logic_scheduler_eusFree_0 & ((! DispatchPlugin_logic_scheduler_arbiters_0_doIt) ? 1'b1 : (~ DispatchPlugin_logic_scheduler_arbiters_0_eusOh)));
  assign DispatchPlugin_logic_scheduler_hartFree_1 = (DispatchPlugin_logic_scheduler_hartFree_0 & (((! DispatchPlugin_logic_candidates_0_ctx_valid) || DispatchPlugin_logic_scheduler_arbiters_0_doIt) ? 1'b1 : (~ 1'b1)));
  assign DispatchPlugin_logic_candidates_0_fire = ((DispatchPlugin_logic_scheduler_arbiters_0_doIt && (! execute_freeze_valid)) && (! DispatchPlugin_api_haltDispatch));
  assign DispatchPlugin_logic_inserter_0_oh = (DispatchPlugin_logic_scheduler_arbiters_0_doIt && DispatchPlugin_logic_scheduler_arbiters_0_eusOh[0]);
  assign DispatchPlugin_logic_inserter_0_trap = DispatchPlugin_logic_candidates_0_ctx_hm_TRAP;
  assign execute_ctrl0_up_LANE_SEL_lane0 = (((|DispatchPlugin_logic_inserter_0_oh) && (! DispatchPlugin_logic_candidates_0_cancel)) && (! DispatchPlugin_api_haltDispatch));
  assign execute_ctrl0_up_Decode_UOP_lane0 = DispatchPlugin_logic_candidates_0_ctx_uop;
  assign execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED;
  assign execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_JUMPED_PC;
  assign execute_ctrl0_up_Prediction_ALIGNED_SLICES_TAKEN_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_TAKEN;
  assign execute_ctrl0_up_Prediction_ALIGNED_SLICES_BRANCH_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_ALIGNED_SLICES_BRANCH;
  assign execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0 = DispatchPlugin_logic_candidates_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0;
  assign execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Prediction_BRANCH_HISTORY;
  assign execute_ctrl0_up_DispatchPlugin_FENCE_OLDER_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_FENCE_OLDER;
  always @(*) begin
    execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_MAY_FLUSH;
    if(when_DispatchPlugin_l439) begin
      execute_ctrl0_up_DispatchPlugin_MAY_FLUSH_lane0 = 1'b0;
    end
  end

  assign execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH;
  assign execute_ctrl0_up_DispatchPlugin_DONT_FLUSH_FROM_LANES_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_DONT_FLUSH_FROM_LANES;
  assign execute_ctrl0_up_DONT_FLUSH_PRECISE_3_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_3;
  assign execute_ctrl0_up_DONT_FLUSH_PRECISE_4_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DONT_FLUSH_PRECISE_4;
  assign execute_ctrl0_up_PC_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_PC;
  assign execute_ctrl0_up_TRAP_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_TRAP;
  assign execute_ctrl0_up_Decode_UOP_ID_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_Decode_UOP_ID;
  assign execute_ctrl0_up_RS1_ENABLE_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RS1_ENABLE;
  assign execute_ctrl0_up_RS1_PHYS_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RS1_PHYS;
  assign execute_ctrl0_up_RS2_ENABLE_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RS2_ENABLE;
  assign execute_ctrl0_up_RS2_PHYS_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RS2_PHYS;
  always @(*) begin
    execute_ctrl0_up_RD_ENABLE_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RD_ENABLE;
    if(when_DispatchPlugin_l439) begin
      execute_ctrl0_up_RD_ENABLE_lane0 = 1'b0;
    end
  end

  assign execute_ctrl0_up_RD_PHYS_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_RD_PHYS;
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0;
  assign execute_ctrl0_up_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_lane0 = DispatchPlugin_logic_candidates_0_ctx_hm_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0;
  assign when_DispatchPlugin_l439 = ((! execute_ctrl0_up_LANE_SEL_lane0) || DispatchPlugin_logic_inserter_0_trap);
  assign execute_ctrl0_up_COMPLETED_lane0 = DispatchPlugin_logic_inserter_0_trap;
  assign DispatchPlugin_logic_inserter_0_layerOhUnfiltred = (DispatchPlugin_logic_inserter_0_oh[0] ? DispatchPlugin_logic_scheduler_arbiters_0_layerOh : 1'b0);
  assign DispatchPlugin_logic_inserter_0_layer_0_1 = DispatchPlugin_logic_inserter_0_layerOhUnfiltred[0];
  assign DispatchPlugin_logic_events_frontendStall = (DispatchPlugin_logic_candidates_0_ctx_valid == 1'b0);
  assign DispatchPlugin_logic_events_backendStall = ((|DispatchPlugin_logic_candidates_0_ctx_valid) && (DispatchPlugin_logic_candidates_0_fire == 1'b0));
  assign _zz_CsrRamPlugin_csrMapper_ramAddress = CsrAccessPlugin_bus_decode_address;
  assign CsrRamPlugin_csrMapper_ramAddress = {(|((_zz_CsrRamPlugin_csrMapper_ramAddress & 12'ha00) == 12'h200)),{(|((_zz_CsrRamPlugin_csrMapper_ramAddress & _zz_CsrRamPlugin_csrMapper_ramAddress_1) == 12'h0)),{(|{_zz_CsrRamPlugin_csrMapper_ramAddress_2,_zz_CsrRamPlugin_csrMapper_ramAddress_3}),(|{_zz_CsrRamPlugin_csrMapper_ramAddress_4,_zz_CsrRamPlugin_csrMapper_ramAddress_5})}}};
  always @(*) begin
    CsrRamPlugin_csrMapper_withRead = 1'b0;
    if(when_CsrAccessPlugin_l252) begin
      CsrRamPlugin_csrMapper_withRead = 1'b1;
    end
  end

  assign CsrRamPlugin_csrMapper_read_valid = (CsrRamPlugin_csrMapper_withRead && (! CsrRamPlugin_api_holdRead));
  assign CsrRamPlugin_csrMapper_read_address = CsrRamPlugin_csrMapper_ramAddress;
  assign when_CsrRamPlugin_l85 = (CsrRamPlugin_csrMapper_withRead && (! CsrRamPlugin_csrMapper_read_ready));
  always @(*) begin
    CsrRamPlugin_csrMapper_doWrite = 1'b0;
    if(when_CsrAccessPlugin_l343_2) begin
      CsrRamPlugin_csrMapper_doWrite = 1'b1;
    end
  end

  assign when_CsrRamPlugin_l92 = (CsrRamPlugin_csrMapper_write_valid && CsrRamPlugin_csrMapper_write_ready);
  assign CsrRamPlugin_csrMapper_write_valid = ((CsrRamPlugin_csrMapper_doWrite && (! CsrRamPlugin_csrMapper_fired)) && (! CsrRamPlugin_api_holdWrite));
  assign CsrRamPlugin_csrMapper_write_address = CsrRamPlugin_csrMapper_ramAddress;
  assign CsrRamPlugin_csrMapper_write_data = CsrAccessPlugin_bus_write_bits;
  assign when_CsrRamPlugin_l96 = ((CsrRamPlugin_csrMapper_doWrite && (! CsrRamPlugin_csrMapper_fired)) && (! CsrRamPlugin_csrMapper_write_ready));
  assign _zz_GSharePlugin_logic_onLearn_hash = LearnPlugin_logic_learn_payload_pcOnLastSlice[15 : 2];
  assign GSharePlugin_logic_onLearn_hash = ({_zz_GSharePlugin_logic_onLearn_hash[0],{_zz_GSharePlugin_logic_onLearn_hash[1],{_zz_GSharePlugin_logic_onLearn_hash[2],{_zz_GSharePlugin_logic_onLearn_hash[3],{_zz_GSharePlugin_logic_onLearn_hash[4],{_zz_GSharePlugin_logic_onLearn_hash[5],{_zz_GSharePlugin_logic_onLearn_hash_1,{_zz_GSharePlugin_logic_onLearn_hash_2,_zz_GSharePlugin_logic_onLearn_hash_3}}}}}}}} ^ _zz_GSharePlugin_logic_onLearn_hash_4);
  assign GSharePlugin_logic_onLearn_incrValue = (LearnPlugin_logic_learn_payload_taken ? 2'b01 : 2'b11);
  always @(*) begin
    GSharePlugin_logic_onLearn_overflow = 1'b0;
    if(when_GSharePlugin_l107) begin
      GSharePlugin_logic_onLearn_overflow = 1'b1;
    end
  end

  assign GSharePlugin_logic_onLearn_updated_0 = (LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 + (1'b1 ? GSharePlugin_logic_onLearn_incrValue : 2'b00));
  assign when_GSharePlugin_l107 = (((LearnPlugin_logic_learn_payload_taken && LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1]) && (! GSharePlugin_logic_onLearn_updated_0[1])) || (((! LearnPlugin_logic_learn_payload_taken) && (! LearnPlugin_logic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0[1])) && GSharePlugin_logic_onLearn_updated_0[1]));
  assign GSharePlugin_logic_mem_write_valid = ((LearnPlugin_logic_learn_valid && LearnPlugin_logic_learn_payload_isBranch) && (! GSharePlugin_logic_onLearn_overflow));
  assign GSharePlugin_logic_mem_write_payload_address = GSharePlugin_logic_onLearn_hash;
  assign GSharePlugin_logic_mem_write_payload_data_0 = GSharePlugin_logic_onLearn_updated_0;
  assign BtbPlugin_logic_onLearn_hash = LearnPlugin_logic_learn_payload_pcOnLastSlice[26 : 11];
  always @(*) begin
    BtbPlugin_logic_memWrite_valid = (LearnPlugin_logic_learn_valid && (LearnPlugin_logic_learn_payload_badPredictedTarget && LearnPlugin_logic_learn_payload_taken));
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_valid = DecoderPlugin_logic_forgetPort_valid;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_address = _zz_BtbPlugin_logic_memWrite_payload_address[8:0];
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_address = _zz_BtbPlugin_logic_memWrite_payload_address_1[8:0];
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_mask = 1'b1;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_mask = 1'b1;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_hash = BtbPlugin_logic_onLearn_hash;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_hash = (~ BtbPlugin_logic_onForget_hash);
    end
  end

  assign BtbPlugin_logic_memWrite_payload_data_0_pcTarget = (LearnPlugin_logic_learn_payload_pcTarget >>> 2'd2);
  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_isBranch = LearnPlugin_logic_learn_payload_isBranch;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_isBranch = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_isPush = LearnPlugin_logic_learn_payload_isPush;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_isPush = 1'b0;
    end
  end

  always @(*) begin
    BtbPlugin_logic_memWrite_payload_data_0_isPop = LearnPlugin_logic_learn_payload_isPop;
    if(DecoderPlugin_logic_forgetPort_valid) begin
      BtbPlugin_logic_memWrite_payload_data_0_isPop = 1'b0;
    end
  end

  assign lane0_integer_WriteBackPlugin_logic_stages_0_hits = {lane0_IntFormatPlugin_logic_stages_0_wb_valid,early0_BranchPlugin_logic_wb_valid};
  assign lane0_integer_WriteBackPlugin_logic_stages_0_muxed = ((lane0_integer_WriteBackPlugin_logic_stages_0_hits[0] ? early0_BranchPlugin_logic_wb_payload : 32'h0) | (lane0_integer_WriteBackPlugin_logic_stages_0_hits[1] ? lane0_IntFormatPlugin_logic_stages_0_wb_payload : 32'h0));
  assign execute_ctrl2_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_valid = (((((execute_ctrl2_down_LANE_SEL_lane0 && execute_ctrl2_down_isReady) && (! execute_lane0_ctrls_2_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_0_hits)) && execute_ctrl2_up_RD_ENABLE_lane0) && execute_ctrl2_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_0_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_hits = lane0_IntFormatPlugin_logic_stages_2_wb_valid;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_muxed = (lane0_integer_WriteBackPlugin_logic_stages_1_hits[0] ? lane0_IntFormatPlugin_logic_stages_2_wb_payload : 32'h0);
  assign lane0_integer_WriteBackPlugin_logic_stages_1_merged = (execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 | lane0_integer_WriteBackPlugin_logic_stages_1_muxed);
  assign execute_ctrl3_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_1_merged;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_valid = (((((execute_ctrl3_down_LANE_SEL_lane0 && execute_ctrl3_down_isReady) && (! execute_lane0_ctrls_3_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_1_hits)) && execute_ctrl3_up_RD_ENABLE_lane0) && execute_ctrl3_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_1_muxed;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_hits = {lane0_IntFormatPlugin_logic_stages_1_wb_valid,CfuPlugin_logic_wb_valid};
  assign lane0_integer_WriteBackPlugin_logic_stages_2_muxed = ((lane0_integer_WriteBackPlugin_logic_stages_2_hits[0] ? CfuPlugin_logic_wb_payload : 32'h0) | (lane0_integer_WriteBackPlugin_logic_stages_2_hits[1] ? lane0_IntFormatPlugin_logic_stages_1_wb_payload : 32'h0));
  assign lane0_integer_WriteBackPlugin_logic_stages_2_merged = (execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 | lane0_integer_WriteBackPlugin_logic_stages_2_muxed);
  assign execute_ctrl4_lane0_integer_WriteBackPlugin_logic_DATA_lane0_bypass = lane0_integer_WriteBackPlugin_logic_stages_2_merged;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_valid = (((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && (|lane0_integer_WriteBackPlugin_logic_stages_2_hits)) && execute_ctrl4_up_RD_ENABLE_lane0) && execute_ctrl4_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data = lane0_integer_WriteBackPlugin_logic_stages_2_muxed;
  assign lane0_integer_WriteBackPlugin_logic_write_port_valid = (((((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_upIsCancel)) && execute_ctrl4_up_RD_ENABLE_lane0) && execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0) && execute_ctrl4_down_COMMIT_lane0);
  assign lane0_integer_WriteBackPlugin_logic_write_port_address = execute_ctrl4_down_RD_PHYS_lane0;
  assign lane0_integer_WriteBackPlugin_logic_write_port_data = execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  assign lane0_integer_WriteBackPlugin_logic_write_port_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign decode_ctrls_1_down_CfuPlugin_logic_CFU_ENABLE_0 = _zz_decode_ctrls_1_down_CfuPlugin_logic_CFU_ENABLE_0[0];
  assign decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_FPU_0[0];
  assign decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0 = _zz_decode_ctrls_1_down_DecoderPlugin_logic_NEED_RM_0[0];
  assign _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h0) == 32'h0);
  assign decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_LANES_LAYER_HIT_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_MAY_FLUSH_0_1[0];
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_1 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00002050) == 32'h00002050);
  assign _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_2 = ((decode_ctrls_1_down_Decode_INSTRUCTION_0 & 32'h00001050) == 32'h00001050);
  assign decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0 = _zz_decode_ctrls_1_down_DispatchPlugin_DONT_FLUSH_FROM_LANES_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0 = _zz_decode_ctrls_1_down_DispatchPlugin_FENCE_OLDER_0[0];
  assign decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_3_0[0];
  assign decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0 = _zz_decode_ctrls_1_down_DONT_FLUSH_PRECISE_4_0_3[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_0_ENABLES_0_0[0];
  assign decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0 = _zz_decode_ctrls_1_down_DispatchPlugin_logic_hcs_0_onRs_1_ENABLES_0_0_1[0];
  assign when_CtrlLaneApi_l50_2 = (decode_ctrls_1_up_isReady || decode_ctrls_1_lane0_upIsCancel);
  assign WhiteboxerPlugin_logic_serializeds_0_fire = (decode_ctrls_1_up_LANE_SEL_0 && (! decode_ctrls_1_up_LANE_SEL_0_regNext_1));
  assign WhiteboxerPlugin_logic_serializeds_0_decodeId = decode_ctrls_1_down_Decode_DOP_ID_0;
  assign WhiteboxerPlugin_logic_serializeds_0_microOpId = decode_ctrls_1_down_Decode_UOP_ID_0;
  assign WhiteboxerPlugin_logic_serializeds_0_microOp = decode_ctrls_1_down_Decode_UOP_0;
  assign when_CtrlLaneApi_l50_3 = (execute_ctrl0_down_isReady || execute_lane0_ctrls_0_downIsCancel);
  assign WhiteboxerPlugin_logic_dispatches_0_fire = (execute_ctrl0_down_LANE_SEL_lane0 && (! execute_ctrl0_down_LANE_SEL_lane0_regNext));
  assign WhiteboxerPlugin_logic_dispatches_0_microOpId = execute_ctrl0_down_Decode_UOP_ID_lane0;
  assign when_CtrlLaneApi_l50_4 = (execute_ctrl2_down_isReady || execute_lane0_ctrls_2_downIsCancel);
  assign WhiteboxerPlugin_logic_executes_0_fire = ((execute_ctrl2_down_LANE_SEL_lane0 && (! execute_ctrl2_down_LANE_SEL_lane0_regNext)) && execute_ctrl2_down_COMMIT_lane0);
  assign WhiteboxerPlugin_logic_executes_0_microOpId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign BtbPlugin_logic_onForget_hash = DecoderPlugin_logic_forgetPort_payload_pcOnLastSlice[26 : 11];
  assign BtbPlugin_logic_memRead_cmd_valid = fetch_logic_ctrls_0_down_isReady;
  assign BtbPlugin_logic_memRead_cmd_payload = _zz_BtbPlugin_logic_memRead_cmd_payload[8:0];
  assign fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS = ((BtbPlugin_logic_memWrite_valid && (BtbPlugin_logic_memWrite_payload_address == BtbPlugin_logic_memRead_cmd_payload)) ? BtbPlugin_logic_memWrite_payload_mask : 1'b0);
  assign fetch_logic_ctrls_0_haltRequest_BtbPlugin_l200 = BtbPlugin_logic_memWrite_valid;
  assign BtbPlugin_logic_predictions = fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0[1];
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash = BtbPlugin_logic_memRead_rsp_0_hash;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget = BtbPlugin_logic_memRead_rsp_0_pcTarget;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch = BtbPlugin_logic_memRead_rsp_0_isBranch;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush = BtbPlugin_logic_memRead_rsp_0_isPush;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop = BtbPlugin_logic_memRead_rsp_0_isPop;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash == fetch_logic_ctrls_1_down_Fetch_WORD_PC[26 : 11]) && 1'b1);
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN = ((! fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) || BtbPlugin_logic_predictions[0]);
  assign BtbPlugin_logic_ras_readIt = fetch_logic_ctrls_0_down_isReady;
  assign BtbPlugin_logic_applyIt_chunksMask = (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && 1'b1);
  assign BtbPlugin_logic_applyIt_chunksTakenOh = (fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN & BtbPlugin_logic_applyIt_chunksMask);
  assign BtbPlugin_logic_applyIt_needIt = (fetch_logic_ctrls_1_up_isValid && (|BtbPlugin_logic_applyIt_chunksTakenOh));
  assign when_BtbPlugin_l233 = (fetch_logic_ctrls_1_up_isReady || fetch_logic_ctrls_1_up_isCancel);
  assign BtbPlugin_logic_applyIt_doIt = (BtbPlugin_logic_applyIt_needIt && (! BtbPlugin_logic_applyIt_correctionSent));
  assign BtbPlugin_logic_applyIt_entry_hash = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_hash;
  assign BtbPlugin_logic_applyIt_entry_pcTarget = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_pcTarget;
  assign BtbPlugin_logic_applyIt_entry_isBranch = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch;
  assign BtbPlugin_logic_applyIt_entry_isPush = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPush;
  assign BtbPlugin_logic_applyIt_entry_isPop = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isPop;
  always @(*) begin
    BtbPlugin_logic_applyIt_pcTarget = BtbPlugin_logic_applyIt_entry_pcTarget;
    if(BtbPlugin_logic_applyIt_entry_isPop) begin
      BtbPlugin_logic_applyIt_pcTarget = BtbPlugin_logic_ras_read;
    end
  end

  assign BtbPlugin_logic_applyIt_rasLogic_pushValid = (BtbPlugin_logic_applyIt_doIt && BtbPlugin_logic_applyIt_entry_isPush);
  assign BtbPlugin_logic_applyIt_rasLogic_pushPc = fetch_logic_ctrls_1_down_Fetch_WORD_PC;
  assign when_BtbPlugin_l246 = (BtbPlugin_logic_applyIt_doIt && BtbPlugin_logic_applyIt_entry_isPop);
  assign BtbPlugin_logic_flushPort_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_logic_flushPort_payload_self = 1'b0;
  assign BtbPlugin_logic_pcPort_valid = BtbPlugin_logic_applyIt_doIt;
  assign BtbPlugin_logic_pcPort_payload_fault = 1'b0;
  assign BtbPlugin_logic_pcPort_payload_pc = ({2'd0,BtbPlugin_logic_applyIt_pcTarget} <<< 2'd2);
  assign fetch_logic_ctrls_1_down_Prediction_WORD_JUMPED = BtbPlugin_logic_applyIt_needIt;
  assign fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_PC = ({2'd0,BtbPlugin_logic_applyIt_pcTarget} <<< 2'd2);
  assign BtbPlugin_logic_applyIt_history_layers_0_history = fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
  assign BtbPlugin_logic_applyIt_history_layersLogic_0_doIt = (BtbPlugin_logic_applyIt_chunksMask[0] && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch);
  assign BtbPlugin_logic_applyIt_history_layersLogic_0_shifted = {BtbPlugin_logic_applyIt_history_layers_0_history[10 : 0],fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN};
  assign BtbPlugin_logic_applyIt_history_layers_1_history = (BtbPlugin_logic_applyIt_history_layersLogic_0_doIt ? BtbPlugin_logic_applyIt_history_layersLogic_0_shifted : BtbPlugin_logic_applyIt_history_layers_0_history);
  assign BtbPlugin_logic_historyPort_valid = ((fetch_logic_ctrls_1_up_isValid && (! BtbPlugin_logic_applyIt_correctionSent)) && (|fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT));
  assign BtbPlugin_logic_historyPort_payload_history = BtbPlugin_logic_applyIt_history_layers_1_history;
  assign fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH[0] = ((fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_hitCalc_HIT && fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_readRsp_ENTRY_isBranch) && 1'b1);
  assign fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN[0] = fetch_logic_ctrls_1_down_BtbPlugin_logic_chunksLogic_0_predict_TAKEN;
  assign AlignerPlugin_logic_nobuffer_flushIt = (|{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign when_AlignerPlugin_l298 = ((AlignerPlugin_logic_nobuffer_flushIt || (! fetch_logic_ctrls_2_down_isValid)) || fetch_logic_ctrls_2_down_isReady);
  assign AlignerPlugin_logic_slices_data_0 = fetch_logic_ctrls_2_down_Fetch_WORD[31 : 0];
  assign AlignerPlugin_logic_slices_mask = ((fetch_logic_ctrls_2_down_valid ? fetch_logic_ctrls_2_down_AlignerPlugin_logic_FETCH_MASK : 1'b0) & 1'b1);
  assign AlignerPlugin_logic_slices_last = 1'b0;
  assign fetch_logic_ctrls_2_down_ready = ((! fetch_logic_ctrls_2_down_valid) || ((decode_ctrls_0_up_isReady && (! AlignerPlugin_api_haltIt)) && (AlignerPlugin_logic_nobuffer_remaningMask == 1'b0)));
  assign AlignerPlugin_logic_extractors_0_ctx_instruction = AlignerPlugin_logic_slicesInstructions_0;
  assign AlignerPlugin_logic_extractors_0_ctx_pc = fetch_logic_ctrls_2_down_Fetch_WORD_PC;
  assign AlignerPlugin_logic_extractors_0_ctx_trap = fetch_logic_ctrls_2_down_TRAP;
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Fetch_ID = fetch_logic_ctrls_2_down_Fetch_ID;
  assign AlignerPlugin_logic_extractors_0_ctx_hm_GSharePlugin_GSHARE_COUNTER_0 = fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0;
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_BRANCH_HISTORY = fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY;
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_BRANCH = fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH;
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_SLICES_TAKEN = fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN;
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMP_PC = fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC;
  assign AlignerPlugin_logic_extractors_0_ctx_hm_Prediction_WORD_JUMPED = fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED;
  assign AlignerPlugin_api_downMoving = decode_ctrls_0_up_isMoving;
  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_read_address = 4'bxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_address = _zz_TrapPlugin_logic_harts_0_crsPorts_read_address;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_read_address = _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign decode_logic_flushes_0_onLanes_0_doIt = (|{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign decode_ctrls_0_lane0_downIsCancel = 1'b0;
  assign decode_ctrls_0_lane0_upIsCancel = decode_logic_flushes_0_onLanes_0_doIt;
  assign decode_logic_flushes_1_onLanes_0_doIt = (|{((DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1) && (1'b0 || (1'b1 && DecoderPlugin_logic_laneLogic_0_flushPort_payload_self))),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign decode_ctrls_1_lane0_downIsCancel = 1'b0;
  assign decode_ctrls_1_lane0_upIsCancel = decode_logic_flushes_1_onLanes_0_doIt;
  assign decode_logic_trapPending[0] = (|{((decode_ctrls_1_up_LANE_SEL_0 && 1'b1) && decode_ctrls_1_down_TRAP_0),((decode_ctrls_0_up_LANE_SEL_0 && 1'b1) && decode_ctrls_0_down_TRAP_0)});
  always @(*) begin
    LsuL1Plugin_logic_banksWrite_address = 9'bxxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_address = {LsuL1Plugin_logic_refill_read_rspAddress[11 : 6],LsuL1Plugin_logic_refill_read_wordIndex};
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 3];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_writeData = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_writeData = LsuL1Plugin_logic_bus_read_rsp_payload_data;
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_writeData[31 : 0] = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
      LsuL1Plugin_logic_banksWrite_writeData[63 : 32] = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_writeMask = 8'bxxxxxxxx;
    LsuL1Plugin_logic_banksWrite_writeMask = 8'hff;
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      LsuL1Plugin_logic_banksWrite_writeMask = 8'h0;
      if(_zz_54[0]) begin
        LsuL1Plugin_logic_banksWrite_writeMask[3 : 0] = execute_ctrl4_down_LsuL1_MASK_lane0;
      end
      if(_zz_54[1]) begin
        LsuL1Plugin_logic_banksWrite_writeMask[7 : 4] = execute_ctrl4_down_LsuL1_MASK_lane0;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
        LsuL1Plugin_logic_banksWrite_writeMask = 8'h0;
      end
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_mask = 4'b0000;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_mask[LsuL1Plugin_logic_refill_read_way] = 1'b1;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_mask = LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      if(LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win) begin
        LsuL1Plugin_logic_waysWrite_mask = 4'b0000;
      end
    end
    if(when_LsuL1Plugin_l1219) begin
      LsuL1Plugin_logic_waysWrite_mask = 4'b1111;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_address = 6'bxxxxxx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_address = LsuL1Plugin_logic_refill_read_rspAddress[11 : 6];
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_address = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
    end
    if(when_LsuL1Plugin_l1219) begin
      LsuL1Plugin_logic_waysWrite_address = LsuL1Plugin_logic_initializer_counter[5:0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_loaded = 1'bx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b1;
    end
    if(when_LsuL1Plugin_l1219) begin
      LsuL1Plugin_logic_waysWrite_tag_loaded = 1'b0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_tag_address = LsuL1Plugin_logic_refill_read_rspAddress[31 : 12];
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_address = _zz_LsuL1Plugin_logic_waysWrite_tag_address;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_waysWrite_tag_fault = 1'bx;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_waysWrite_tag_fault = LsuL1Plugin_logic_refill_read_faulty;
      end
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_waysWrite_tag_fault = _zz_LsuL1Plugin_logic_waysWrite_tag_fault;
    end
  end

  assign LsuL1Plugin_logic_waysWrite_valid = (|LsuL1Plugin_logic_waysWrite_mask);
  assign LsuL1Plugin_logic_banks_0_write_valid = LsuL1Plugin_logic_banksWrite_mask[0];
  assign LsuL1Plugin_logic_banks_0_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_0_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_0_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_0_read_rsp = LsuL1Plugin_logic_banks_0_mem_rd_data;
  assign LsuL1Plugin_logic_banks_1_write_valid = LsuL1Plugin_logic_banksWrite_mask[1];
  assign LsuL1Plugin_logic_banks_1_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_1_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_1_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_1_read_rsp = LsuL1Plugin_logic_banks_1_mem_rd_data;
  assign LsuL1Plugin_logic_banks_2_write_valid = LsuL1Plugin_logic_banksWrite_mask[2];
  assign LsuL1Plugin_logic_banks_2_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_2_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_2_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_2_read_rsp = LsuL1Plugin_logic_banks_2_mem_rd_data;
  assign LsuL1Plugin_logic_banks_3_write_valid = LsuL1Plugin_logic_banksWrite_mask[3];
  assign LsuL1Plugin_logic_banks_3_write_payload_address = LsuL1Plugin_logic_banksWrite_address;
  assign LsuL1Plugin_logic_banks_3_write_payload_data = LsuL1Plugin_logic_banksWrite_writeData;
  assign LsuL1Plugin_logic_banks_3_write_payload_mask = LsuL1Plugin_logic_banksWrite_writeMask;
  assign LsuL1Plugin_logic_banks_3_read_rsp = LsuL1Plugin_logic_banks_3_mem_rd_data;
  assign _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_0_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_1_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_ways_2_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_2_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_2_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_2_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_2_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_2_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_2_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_2_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_ways_3_lsuRead_rsp_loaded = LsuL1Plugin_logic_ways_3_mem_spinal_port1;
  assign LsuL1Plugin_logic_ways_3_lsuRead_rsp_loaded = _zz_LsuL1Plugin_logic_ways_3_lsuRead_rsp_loaded[0];
  assign LsuL1Plugin_logic_ways_3_lsuRead_rsp_address = _zz_LsuL1Plugin_logic_ways_3_lsuRead_rsp_loaded[20 : 1];
  assign LsuL1Plugin_logic_ways_3_lsuRead_rsp_fault = _zz_LsuL1Plugin_logic_ways_3_lsuRead_rsp_loaded[21];
  assign _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_dirty = LsuL1Plugin_logic_shared_mem_spinal_port1;
  assign _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_dirty[2 : 0];
  assign LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0 = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0[0 : 0];
  assign LsuL1Plugin_logic_shared_lsuRead_rsp_plru_1 = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0[2 : 1];
  assign LsuL1Plugin_logic_shared_lsuRead_rsp_dirty = _zz_LsuL1Plugin_logic_shared_lsuRead_rsp_dirty[6 : 3];
  always @(*) begin
    LsuL1Plugin_logic_refill_slots_0_loadedSet = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_refill_slots_0_loadedSet = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_refill_slots_0_loadedDone = (LsuL1Plugin_logic_refill_slots_0_loadedCounter == 1'b1);
  assign LsuL1Plugin_logic_refill_slots_0_free = ((! LsuL1Plugin_logic_refill_slots_0_valid) && 1'b1);
  assign LsuL1Plugin_logic_refill_slots_0_fire = ((! execute_freeze_valid) && LsuL1Plugin_logic_refill_slots_0_loadedDone);
  assign LsuL1Plugin_logic_refill_free = LsuL1Plugin_logic_refill_slots_0_free;
  assign LsuL1Plugin_logic_refill_full = (&(! LsuL1Plugin_logic_refill_slots_0_free));
  assign when_LsuL1Plugin_l377 = (LsuL1Plugin_logic_refill_push_valid && LsuL1Plugin_logic_refill_free[0]);
  assign when_LsuL1Plugin_l381 = LsuL1Plugin_logic_refill_free[0];
  assign LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0 = ((LsuL1Plugin_logic_refill_slots_0_valid && (! LsuL1Plugin_logic_refill_slots_0_cmdSent)) && (LsuL1Plugin_logic_refill_slots_0_victim == 1'b0));
  assign LsuL1Plugin_logic_refill_read_arbiter_hits = LsuL1Plugin_logic_refill_read_arbiter_slotsWithId_0_0;
  assign LsuL1Plugin_logic_refill_read_arbiter_hit = (|LsuL1Plugin_logic_refill_read_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_refill_read_arbiter_oh = (LsuL1Plugin_logic_refill_read_arbiter_hits & 1'b1);
    if(when_LsuL1Plugin_l301) begin
      LsuL1Plugin_logic_refill_read_arbiter_oh = LsuL1Plugin_logic_refill_read_arbiter_lock;
    end
  end

  assign when_LsuL1Plugin_l301 = (|LsuL1Plugin_logic_refill_read_arbiter_lock);
  assign LsuL1Plugin_logic_bus_read_cmd_fire = (LsuL1Plugin_logic_bus_read_cmd_valid && LsuL1Plugin_logic_bus_read_cmd_ready);
  assign LsuL1Plugin_logic_refill_read_cmdAddress = {LsuL1Plugin_logic_refill_slots_0_address[31 : 6],6'h0};
  assign LsuL1Plugin_logic_bus_read_cmd_valid = LsuL1Plugin_logic_refill_read_arbiter_hit;
  assign LsuL1Plugin_logic_bus_read_cmd_payload_address = LsuL1Plugin_logic_refill_read_cmdAddress;
  assign LsuL1Plugin_logic_refill_read_rspAddress = LsuL1Plugin_logic_refill_slots_0_address;
  assign LsuL1Plugin_logic_refill_read_dirty = LsuL1Plugin_logic_refill_slots_0_dirty;
  assign LsuL1Plugin_logic_refill_read_way = LsuL1Plugin_logic_refill_slots_0_way;
  assign LsuL1Plugin_logic_refill_read_rspWithData = 1'b1;
  always @(*) begin
    LsuL1Plugin_logic_refill_read_writeReservation_take = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      LsuL1Plugin_logic_refill_read_writeReservation_take = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_read_bankWriteNotif[0] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 2'b00));
    LsuL1Plugin_logic_refill_read_bankWriteNotif[1] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 2'b01));
    LsuL1Plugin_logic_refill_read_bankWriteNotif[2] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 2'b10));
    LsuL1Plugin_logic_refill_read_bankWriteNotif[3] = ((LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_refill_read_rspWithData) && (LsuL1Plugin_logic_refill_read_way == 2'b11));
  end

  always @(*) begin
    LsuL1Plugin_logic_banksWrite_mask[0] = LsuL1Plugin_logic_refill_read_bankWriteNotif[0];
    LsuL1Plugin_logic_banksWrite_mask[1] = LsuL1Plugin_logic_refill_read_bankWriteNotif[1];
    LsuL1Plugin_logic_banksWrite_mask[2] = LsuL1Plugin_logic_refill_read_bankWriteNotif[2];
    LsuL1Plugin_logic_banksWrite_mask[3] = LsuL1Plugin_logic_refill_read_bankWriteNotif[3];
    if(LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win) begin
      if(when_LsuL1Plugin_l929) begin
        LsuL1Plugin_logic_banksWrite_mask[0] = ((2'b00 == LsuL1Plugin_logic_lsu_ctrl_wayId) && LsuL1Plugin_logic_lsu_ctrl_doWrite);
      end
      if(when_LsuL1Plugin_l929_1) begin
        LsuL1Plugin_logic_banksWrite_mask[1] = ((2'b01 == LsuL1Plugin_logic_lsu_ctrl_wayId) && LsuL1Plugin_logic_lsu_ctrl_doWrite);
      end
      if(when_LsuL1Plugin_l929_2) begin
        LsuL1Plugin_logic_banksWrite_mask[2] = ((2'b10 == LsuL1Plugin_logic_lsu_ctrl_wayId) && LsuL1Plugin_logic_lsu_ctrl_doWrite);
      end
      if(when_LsuL1Plugin_l929_3) begin
        LsuL1Plugin_logic_banksWrite_mask[3] = ((2'b11 == LsuL1Plugin_logic_lsu_ctrl_wayId) && LsuL1Plugin_logic_lsu_ctrl_doWrite);
      end
    end
  end

  assign when_LsuL1Plugin_l450 = (LsuL1Plugin_logic_bus_read_rsp_valid && LsuL1Plugin_logic_bus_read_rsp_payload_error);
  always @(*) begin
    LsuL1Plugin_logic_refill_read_fire = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_refill_read_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_read_reservation_take = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_refill_read_reservation_take = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_refill_read_faulty = (LsuL1Plugin_logic_refill_read_hadError || LsuL1Plugin_logic_bus_read_rsp_payload_error);
  always @(*) begin
    LsuL1Plugin_logic_refillCompletions = 1'b0;
    if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
      if(when_LsuL1Plugin_l463) begin
        LsuL1Plugin_logic_refillCompletions[0] = 1'b1;
      end
    end
  end

  assign LsuL1Plugin_logic_bus_read_rsp_ready = 1'b1;
  assign when_LsuL1Plugin_l463 = ((LsuL1Plugin_logic_refill_read_wordIndex == 3'b111) || (! LsuL1Plugin_logic_refill_read_rspWithData));
  assign LsuL1_REFILL_BUSY = ((! LsuL1Plugin_logic_refill_slots_0_loaded) && (! LsuL1Plugin_logic_refill_slots_0_loadedSet));
  always @(*) begin
    LsuL1Plugin_logic_writeback_slots_0_fire = 1'b0;
    if(LsuL1Plugin_logic_bus_write_rsp_valid) begin
      LsuL1Plugin_logic_writeback_slots_0_fire = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_writeback_slots_0_timer_done = (LsuL1Plugin_logic_writeback_slots_0_timer_counter == 1'b1);
  assign when_LsuL1Plugin_l530 = (LsuL1Plugin_logic_writeback_slots_0_timer_done && (LsuL1Plugin_logic_writeback_slots_0_fire || (! LsuL1Plugin_logic_writeback_slots_0_busy)));
  assign LsuL1Plugin_logic_writeback_slots_0_free = (! LsuL1Plugin_logic_writeback_slots_0_valid);
  assign LsuL1_WRITEBACK_BUSY = (LsuL1Plugin_logic_writeback_slots_0_valid || LsuL1Plugin_logic_writeback_slots_0_fire);
  assign LsuL1Plugin_logic_writebackBusy = (|LsuL1Plugin_logic_writeback_slots_0_valid);
  assign LsuL1Plugin_logic_writeback_free = LsuL1Plugin_logic_writeback_slots_0_free;
  assign LsuL1Plugin_logic_writeback_full = (&(! LsuL1Plugin_logic_writeback_slots_0_free));
  always @(*) begin
    LsuL1Plugin_logic_writeback_push_valid = 1'b0;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_valid = LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_writeback_push_valid = 1'b0;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_writeback_push_payload_address = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_payload_address = ({6'd0,{_zz_LsuL1Plugin_logic_waysWrite_tag_address,execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]}} <<< 3'd6);
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_payload_address = ({6'd0,{_zz_LsuL1Plugin_logic_writeback_push_payload_address,execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]}} <<< 3'd6);
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_writeback_push_payload_way = 2'bxx;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_writeback_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_needFlushSel;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_writeback_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_targetWay;
    end
  end

  assign when_LsuL1Plugin_l556 = (LsuL1Plugin_logic_writeback_free[0] && LsuL1Plugin_logic_writeback_push_valid);
  assign when_LsuL1Plugin_l561 = LsuL1Plugin_logic_writeback_free[0];
  assign LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0 = (LsuL1Plugin_logic_writeback_slots_0_valid && (! LsuL1Plugin_logic_writeback_slots_0_readCmdDone));
  assign LsuL1Plugin_logic_writeback_read_arbiter_hits = LsuL1Plugin_logic_writeback_read_arbiter_slotsWithId_0_0;
  assign LsuL1Plugin_logic_writeback_read_arbiter_hit = (|LsuL1Plugin_logic_writeback_read_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_writeback_read_arbiter_oh = (LsuL1Plugin_logic_writeback_read_arbiter_hits & 1'b1);
    if(when_LsuL1Plugin_l301_1) begin
      LsuL1Plugin_logic_writeback_read_arbiter_oh = LsuL1Plugin_logic_writeback_read_arbiter_lock;
    end
  end

  assign when_LsuL1Plugin_l301_1 = (|LsuL1Plugin_logic_writeback_read_arbiter_lock);
  assign LsuL1Plugin_logic_writeback_read_address = LsuL1Plugin_logic_writeback_slots_0_address;
  assign LsuL1Plugin_logic_writeback_read_way = LsuL1Plugin_logic_writeback_slots_0_way;
  assign LsuL1Plugin_logic_writeback_read_slotRead_valid = LsuL1Plugin_logic_writeback_read_arbiter_hit;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex = LsuL1Plugin_logic_writeback_read_wordIndex;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_way = LsuL1Plugin_logic_writeback_read_way;
  assign LsuL1Plugin_logic_writeback_read_slotRead_payload_last = (LsuL1Plugin_logic_writeback_read_wordIndex == 3'b111);
  assign when_LsuL1Plugin_l605 = (LsuL1Plugin_logic_writeback_read_slotRead_valid && LsuL1Plugin_logic_writeback_read_slotRead_payload_last);
  always @(*) begin
    LsuL1Plugin_logic_banks_0_read_cmd_valid = LsuL1Plugin_logic_banks_0_usedByWriteback;
    if(when_LsuL1Plugin_l718) begin
      LsuL1Plugin_logic_banks_0_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_0_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 2'b00));
  always @(*) begin
    LsuL1Plugin_logic_banks_0_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l719) begin
      LsuL1Plugin_logic_banks_0_read_cmd_payload = LsuL1Plugin_logic_lsu_rb0_readAddress;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_1_read_cmd_valid = LsuL1Plugin_logic_banks_1_usedByWriteback;
    if(when_LsuL1Plugin_l718_1) begin
      LsuL1Plugin_logic_banks_1_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_1_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 2'b01));
  always @(*) begin
    LsuL1Plugin_logic_banks_1_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l719_1) begin
      LsuL1Plugin_logic_banks_1_read_cmd_payload = LsuL1Plugin_logic_lsu_rb0_readAddress;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_2_read_cmd_valid = LsuL1Plugin_logic_banks_2_usedByWriteback;
    if(when_LsuL1Plugin_l718_2) begin
      LsuL1Plugin_logic_banks_2_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_2_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 2'b10));
  always @(*) begin
    LsuL1Plugin_logic_banks_2_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l719_2) begin
      LsuL1Plugin_logic_banks_2_read_cmd_payload = LsuL1Plugin_logic_lsu_rb0_readAddress;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_banks_3_read_cmd_valid = LsuL1Plugin_logic_banks_3_usedByWriteback;
    if(when_LsuL1Plugin_l718_3) begin
      LsuL1Plugin_logic_banks_3_read_cmd_valid = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_banks_3_usedByWriteback = (LsuL1Plugin_logic_writeback_read_slotRead_valid && (LsuL1Plugin_logic_writeback_read_way == 2'b11));
  always @(*) begin
    LsuL1Plugin_logic_banks_3_read_cmd_payload = {LsuL1Plugin_logic_writeback_read_address[11 : 6],LsuL1Plugin_logic_writeback_read_wordIndex};
    if(when_LsuL1Plugin_l719_3) begin
      LsuL1Plugin_logic_banks_3_read_cmd_payload = LsuL1Plugin_logic_lsu_rb0_readAddress;
    end
  end

  assign LsuL1Plugin_logic_writeback_read_readedData = _zz_LsuL1Plugin_logic_writeback_read_readedData;
  assign LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0 = ((LsuL1Plugin_logic_writeback_slots_0_valid && LsuL1Plugin_logic_writeback_slots_0_victimBufferReady) && (! LsuL1Plugin_logic_writeback_slots_0_writeCmdDone));
  assign LsuL1Plugin_logic_writeback_write_arbiter_hits = LsuL1Plugin_logic_writeback_write_arbiter_slotsWithId_0_0;
  assign LsuL1Plugin_logic_writeback_write_arbiter_hit = (|LsuL1Plugin_logic_writeback_write_arbiter_hits);
  always @(*) begin
    LsuL1Plugin_logic_writeback_write_arbiter_oh = (LsuL1Plugin_logic_writeback_write_arbiter_hits & 1'b1);
    if(when_LsuL1Plugin_l301_2) begin
      LsuL1Plugin_logic_writeback_write_arbiter_oh = LsuL1Plugin_logic_writeback_write_arbiter_lock;
    end
  end

  assign when_LsuL1Plugin_l301_2 = (|LsuL1Plugin_logic_writeback_write_arbiter_lock);
  assign LsuL1Plugin_logic_writeback_write_last = (LsuL1Plugin_logic_writeback_write_wordIndex == 3'b111);
  assign LsuL1Plugin_logic_writeback_write_bufferRead_valid = LsuL1Plugin_logic_writeback_write_arbiter_hit;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_payload_last = LsuL1Plugin_logic_writeback_write_last;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_payload_address = LsuL1Plugin_logic_writeback_slots_0_address;
  assign LsuL1Plugin_logic_writeback_write_bufferRead_fire = (LsuL1Plugin_logic_writeback_write_bufferRead_valid && LsuL1Plugin_logic_writeback_write_bufferRead_ready);
  assign when_LsuL1Plugin_l676 = (LsuL1Plugin_logic_writeback_write_bufferRead_fire && LsuL1Plugin_logic_writeback_write_last);
  always @(*) begin
    LsuL1Plugin_logic_writeback_write_bufferRead_ready = LsuL1Plugin_logic_writeback_write_cmd_ready;
    if(when_Stream_l399) begin
      LsuL1Plugin_logic_writeback_write_bufferRead_ready = 1'b1;
    end
  end

  assign when_Stream_l399 = (! LsuL1Plugin_logic_writeback_write_cmd_valid);
  assign LsuL1Plugin_logic_writeback_write_cmd_valid = LsuL1Plugin_logic_writeback_write_bufferRead_rValid;
  assign LsuL1Plugin_logic_writeback_write_cmd_payload_address = LsuL1Plugin_logic_writeback_write_bufferRead_rData_address;
  assign LsuL1Plugin_logic_writeback_write_cmd_payload_last = LsuL1Plugin_logic_writeback_write_bufferRead_rData_last;
  assign _zz_LsuL1Plugin_logic_writeback_write_word = LsuL1Plugin_logic_writeback_write_wordIndex;
  assign LsuL1Plugin_logic_writeback_write_word = LsuL1Plugin_logic_writeback_victimBuffer_spinal_port1;
  assign LsuL1Plugin_logic_bus_write_cmd_valid = LsuL1Plugin_logic_writeback_write_cmd_valid;
  assign LsuL1Plugin_logic_writeback_write_cmd_ready = LsuL1Plugin_logic_bus_write_cmd_ready;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address = LsuL1Plugin_logic_writeback_write_cmd_payload_address;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data = LsuL1Plugin_logic_writeback_write_word;
  assign LsuL1Plugin_logic_bus_write_cmd_payload_last = LsuL1Plugin_logic_writeback_write_cmd_payload_last;
  assign LsuL1Plugin_logic_lsu_rb0_readAddress = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 3];
  always @(*) begin
    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[0] = LsuL1Plugin_logic_banks_0_usedByWriteback;
    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[1] = LsuL1Plugin_logic_banks_1_usedByWriteback;
    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[2] = LsuL1Plugin_logic_banks_2_usedByWriteback;
    execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0[3] = LsuL1Plugin_logic_banks_3_usedByWriteback;
  end

  assign when_LsuL1Plugin_l718 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l719 = (! LsuL1Plugin_logic_banks_0_usedByWriteback);
  assign when_LsuL1Plugin_l718_1 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l719_1 = (! LsuL1Plugin_logic_banks_1_usedByWriteback);
  assign when_LsuL1Plugin_l718_2 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l719_2 = (! LsuL1Plugin_logic_banks_2_usedByWriteback);
  assign when_LsuL1Plugin_l718_3 = (! execute_freeze_valid);
  assign when_LsuL1Plugin_l719_3 = (! LsuL1Plugin_logic_banks_3_usedByWriteback);
  assign when_LsuL1Plugin_l735 = (! execute_freeze_valid);
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_0 = LsuL1Plugin_logic_banks_0_read_rsp;
  always @(*) begin
    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[0] = (execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[2'b00] || LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg);
    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[1] = (execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[2'b01] || LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg);
    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[2] = (execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[2'b10] || LsuL1Plugin_logic_lsu_rb1_onBanks_2_busyReg);
    execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0[3] = (execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0[2'b11] || LsuL1Plugin_logic_lsu_rb1_onBanks_3_busyReg);
  end

  assign when_LsuL1Plugin_l735_1 = (! execute_freeze_valid);
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_1 = LsuL1Plugin_logic_banks_1_read_rsp;
  assign when_LsuL1Plugin_l735_2 = (! execute_freeze_valid);
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_2 = LsuL1Plugin_logic_banks_2_read_rsp;
  assign when_LsuL1Plugin_l735_3 = (! execute_freeze_valid);
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_WORDS_lane0_3 = LsuL1Plugin_logic_banks_3_read_rsp;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2 = _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3 = _zz_execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3;
  assign _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0];
  assign _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1];
  assign _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_2 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[2];
  assign _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_3 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[3];
  assign execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 = (((_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0 ? execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 : 32'h0) | (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 ? execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 : 32'h0)) | ((_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_2 ? execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2 : 32'h0) | (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_3 ? execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3 : 32'h0)));
  always @(*) begin
    execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[0] = ((execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 && (execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0[31 : 2] == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 2])) && 1'b1);
    execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[1] = ((execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 && (execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0[31 : 2] == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 2])) && 1'b1);
  end

  assign LsuL1Plugin_logic_shared_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_shared_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0 = (LsuL1Plugin_logic_shared_write_valid && (LsuL1Plugin_logic_shared_write_payload_address == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]));
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 = LsuL1Plugin_logic_shared_write_payload_data_plru_0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_1 = LsuL1Plugin_logic_shared_write_payload_data_plru_1;
  assign execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty = LsuL1Plugin_logic_shared_write_payload_data_dirty;
  assign LsuL1Plugin_logic_ways_0_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_0_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign LsuL1Plugin_logic_ways_1_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_1_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign LsuL1Plugin_logic_ways_2_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_2_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  assign LsuL1Plugin_logic_ways_3_lsuRead_cmd_valid = (! execute_freeze_valid);
  assign LsuL1Plugin_logic_ways_3_lsuRead_cmd_payload = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
  always @(*) begin
    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 = LsuL1Plugin_logic_shared_lsuRead_rsp_plru_0;
    if(execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0) begin
      execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 = execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
    end
  end

  always @(*) begin
    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_1 = LsuL1Plugin_logic_shared_lsuRead_rsp_plru_1;
    if(execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0) begin
      execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_1 = execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_1;
    end
  end

  always @(*) begin
    execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty = LsuL1Plugin_logic_shared_lsuRead_rsp_dirty;
    if(execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0) begin
      execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty = execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
    end
  end

  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded = LsuL1Plugin_logic_ways_0_lsuRead_rsp_loaded;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address = LsuL1Plugin_logic_ways_0_lsuRead_rsp_address;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault = LsuL1Plugin_logic_ways_0_lsuRead_rsp_fault;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded = LsuL1Plugin_logic_ways_1_lsuRead_rsp_loaded;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address = LsuL1Plugin_logic_ways_1_lsuRead_rsp_address;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault = LsuL1Plugin_logic_ways_1_lsuRead_rsp_fault;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded = LsuL1Plugin_logic_ways_2_lsuRead_rsp_loaded;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address = LsuL1Plugin_logic_ways_2_lsuRead_rsp_address;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault = LsuL1Plugin_logic_ways_2_lsuRead_rsp_fault;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded = LsuL1Plugin_logic_ways_3_lsuRead_rsp_loaded;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address = LsuL1Plugin_logic_ways_3_lsuRead_rsp_address;
  assign execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault = LsuL1Plugin_logic_ways_3_lsuRead_rsp_fault;
  assign LsuL1Plugin_logic_lsu_sharedBypassers_0_hit = (LsuL1Plugin_logic_shared_write_valid && (LsuL1Plugin_logic_shared_write_payload_address == execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6]));
  assign execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_0 = (LsuL1Plugin_logic_lsu_sharedBypassers_0_hit ? LsuL1Plugin_logic_shared_write_payload_data_plru_0 : execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_0);
  assign execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_plru_1 = (LsuL1Plugin_logic_lsu_sharedBypassers_0_hit ? LsuL1Plugin_logic_shared_write_payload_data_plru_1 : execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_plru_1);
  assign execute_ctrl3_LsuL1Plugin_logic_SHARED_lane0_bypass_dirty = (LsuL1Plugin_logic_lsu_sharedBypassers_0_hit ? LsuL1Plugin_logic_shared_write_payload_data_dirty : execute_ctrl3_up_LsuL1Plugin_logic_SHARED_lane0_dirty);
  always @(*) begin
    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0] = (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded && (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1] = (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded && (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[2] = (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded && (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
    execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0[3] = (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded && (execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address == execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0[31 : 12]));
  end

  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 = (|execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0);
  assign execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0 = (execute_ctrl4_down_LsuL1_STORE_lane0 || execute_ctrl4_down_LsuL1_ATOMIC_lane0);
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_0_state = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_0[0];
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0 = (! LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_0_state);
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_1_stateSel = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0;
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_1_state = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_1[LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_1_stateSel];
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_1 = (! LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_logic_1_state);
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_evict_id = {LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_0,LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_evict_sel_1};
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_0[0] = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id[1];
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_update_logic_1_sel = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id[1 : 1];
  always @(*) begin
    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_1 = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_1;
    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_1[LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_update_logic_1_sel] = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id[0];
  end

  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_0 = execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  assign LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_context_state_1 = execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_1;
  always @(*) begin
    LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take = 1'b0;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_take = 1'b1;
    end
  end

  assign LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_take = 1'b0;
  assign LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_evict_id;
  assign LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback = _zz_LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback[LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate];
  assign LsuL1Plugin_logic_lsu_ctrl_refillHazards = (LsuL1Plugin_logic_refill_slots_0_valid && (LsuL1Plugin_logic_refill_slots_0_address[11 : 6] == execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6]));
  assign LsuL1Plugin_logic_lsu_ctrl_writebackHazards = (LsuL1Plugin_logic_writeback_slots_0_valid && (LsuL1Plugin_logic_writeback_slots_0_address[11 : 6] == execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[11 : 6]));
  assign LsuL1Plugin_logic_lsu_ctrl_refillHazard = (|LsuL1Plugin_logic_lsu_ctrl_refillHazards);
  assign LsuL1Plugin_logic_lsu_ctrl_writebackHazard = (|LsuL1Plugin_logic_lsu_ctrl_writebackHazards);
  assign LsuL1Plugin_logic_lsu_ctrl_wasDirty = (|(execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty & execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_loadedDirties = ({execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded,{execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded,{execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded,execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded}}} & execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty);
  assign LsuL1Plugin_logic_lsu_ctrl_refillWayWasDirty = LsuL1Plugin_logic_lsu_ctrl_loadedDirties[LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate];
  assign LsuL1Plugin_logic_lsu_ctrl_writeToReadHazard = 1'b0;
  assign LsuL1Plugin_logic_lsu_ctrl_bankNotRead = (|(execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 & execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_loadHazard = ((execute_ctrl4_down_LsuL1_LOAD_lane0 && (! execute_ctrl4_down_LsuL1_PREFETCH_lane0)) && (LsuL1Plugin_logic_lsu_ctrl_bankNotRead || LsuL1Plugin_logic_lsu_ctrl_writeToReadHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_storeHazard = ((execute_ctrl4_down_LsuL1_STORE_lane0 && (! execute_ctrl4_down_LsuL1_PREFETCH_lane0)) && (! LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win));
  assign LsuL1Plugin_logic_lsu_ctrl_preventSideEffects = (execute_ctrl4_down_LsuL1_ABORD_lane0 || execute_freeze_valid);
  assign LsuL1Plugin_logic_lsu_ctrl_flushHazard = (execute_ctrl4_down_LsuL1_FLUSH_lane0 && (! LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win));
  assign LsuL1Plugin_logic_lsu_ctrl_coherencyHazard = 1'b0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0 = 1'b0;
  assign execute_ctrl4_down_LsuL1_HAZARD_lane0 = (((((LsuL1Plugin_logic_lsu_ctrl_hazardReg || LsuL1Plugin_logic_lsu_ctrl_loadHazard) || LsuL1Plugin_logic_lsu_ctrl_refillHazard) || LsuL1Plugin_logic_lsu_ctrl_storeHazard) || LsuL1Plugin_logic_lsu_ctrl_coherencyHazard) || execute_ctrl4_down_LsuL1Plugin_logic_HAZARD_FORCED_lane0);
  assign execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0 = (LsuL1Plugin_logic_lsu_ctrl_flushHazardReg || LsuL1Plugin_logic_lsu_ctrl_flushHazard);
  assign execute_ctrl4_down_LsuL1_MISS_lane0 = (! execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0);
  assign execute_ctrl4_down_LsuL1_FAULT_lane0 = ((execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && (|(execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 & {execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault,{execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault,{execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault,execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault}}}))) && (! execute_ctrl4_down_LsuL1_FLUSH_lane0));
  assign execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0 = ((execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0) && 1'b0);
  assign execute_ctrl4_down_LsuL1_REFILL_HIT_lane0 = LsuL1Plugin_logic_lsu_ctrl_refillHazard;
  assign LsuL1Plugin_logic_events_loadAccess = ((((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_isReady) && (! execute_lane0_ctrls_4_upIsCancel)) && execute_ctrl4_down_LsuL1_SEL_lane0) && execute_ctrl4_down_LsuL1_LOAD_lane0);
  assign LsuL1Plugin_logic_events_loadMiss = ((LsuL1Plugin_logic_events_loadAccess && (! execute_ctrl4_down_LsuL1_HAZARD_lane0)) && execute_ctrl4_down_LsuL1_MISS_lane0);
  assign LsuL1Plugin_logic_lsu_ctrl_canRefill = (((! (LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback && LsuL1Plugin_logic_writeback_full)) && (! LsuL1Plugin_logic_refill_full)) && (! LsuL1Plugin_logic_lsu_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_canFlush = (((LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win && (! LsuL1Plugin_logic_writeback_full)) && (! (|LsuL1Plugin_logic_refill_slots_0_valid))) && (! LsuL1Plugin_logic_lsu_ctrl_writebackHazard));
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs = LsuL1Plugin_logic_lsu_ctrl_loadedDirties;
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0 = LsuL1Plugin_logic_lsu_ctrl_needFlushs;
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0 = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0[0];
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1 = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0[1];
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_2 = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0[2];
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_3 = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0[3];
  always @(*) begin
    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh[0] = (LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0 && (! 1'b0));
    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh[1] = (LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1 && (! LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0));
    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh[2] = (LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_2 && (! LsuL1Plugin_logic_lsu_ctrl_needFlushs_range_0_to_1));
    _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh[3] = (LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_3 && (! LsuL1Plugin_logic_lsu_ctrl_needFlushs_range_0_to_2));
  end

  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_range_0_to_1 = (|{LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1,LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0});
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushs_range_0_to_2 = (|{LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_2,{LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_1,LsuL1Plugin_logic_lsu_ctrl_needFlushs_bools_0}});
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushOh = _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushOh;
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel = LsuL1Plugin_logic_lsu_ctrl_needFlushOh[3];
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel_1 = (LsuL1Plugin_logic_lsu_ctrl_needFlushOh[1] || _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel);
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel_2 = (LsuL1Plugin_logic_lsu_ctrl_needFlushOh[2] || _zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel);
  assign LsuL1Plugin_logic_lsu_ctrl_needFlushSel = {_zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel_2,_zz_LsuL1Plugin_logic_lsu_ctrl_needFlushSel_1};
  assign LsuL1Plugin_logic_lsu_ctrl_isAccess = (((! execute_ctrl4_down_LsuL1_FLUSH_lane0) && (! execute_ctrl4_down_LsuL1_CLEAN_lane0)) && (! execute_ctrl4_down_LsuL1_INVALID_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_askRefill = ((LsuL1Plugin_logic_lsu_ctrl_isAccess && execute_ctrl4_down_LsuL1_MISS_lane0) && LsuL1Plugin_logic_lsu_ctrl_canRefill);
  assign LsuL1Plugin_logic_lsu_ctrl_askUpgrade = ((LsuL1Plugin_logic_lsu_ctrl_isAccess && execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0) && LsuL1Plugin_logic_lsu_ctrl_canRefill);
  assign LsuL1Plugin_logic_lsu_ctrl_askFlush = ((execute_ctrl4_down_LsuL1_FLUSH_lane0 && LsuL1Plugin_logic_lsu_ctrl_canFlush) && (|LsuL1Plugin_logic_lsu_ctrl_needFlushs));
  assign LsuL1Plugin_logic_lsu_ctrl_askCbm = (execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0 && (execute_ctrl4_down_LsuL1_INVALID_lane0 || (execute_ctrl4_down_LsuL1_CLEAN_lane0 && LsuL1Plugin_logic_lsu_ctrl_wasDirty)));
  assign LsuL1Plugin_logic_lsu_ctrl_doRefill = (execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askRefill);
  assign LsuL1Plugin_logic_lsu_ctrl_doUpgrade = (execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askUpgrade);
  assign LsuL1Plugin_logic_lsu_ctrl_doFlush = (execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askFlush);
  assign LsuL1Plugin_logic_lsu_ctrl_doWrite = ((((execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuL1_STORE_lane0) && execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HIT_lane0) && _zz_LsuL1Plugin_logic_lsu_ctrl_doWrite[0]) && (! execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0));
  assign LsuL1Plugin_logic_lsu_ctrl_doCbm = (((((execute_ctrl4_down_LsuL1_SEL_lane0 && LsuL1Plugin_logic_lsu_ctrl_askCbm) && LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win) && (! LsuL1Plugin_logic_writeback_full)) && (! LsuL1Plugin_logic_lsu_ctrl_refillHazard)) && (! LsuL1Plugin_logic_lsu_ctrl_writebackHazard));
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_wayId = (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_1 || _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_3);
  assign _zz_LsuL1Plugin_logic_lsu_ctrl_wayId_1 = (_zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_2 || _zz_execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0_3);
  assign LsuL1Plugin_logic_lsu_ctrl_wayId = {_zz_LsuL1Plugin_logic_lsu_ctrl_wayId_1,_zz_LsuL1Plugin_logic_lsu_ctrl_wayId};
  assign LsuL1Plugin_logic_lsu_ctrl_targetWay = (LsuL1Plugin_logic_lsu_ctrl_askUpgrade ? LsuL1Plugin_logic_lsu_ctrl_wayId : LsuL1Plugin_logic_lsu_ctrl_refillWayWithoutUpdate);
  assign _zz_45 = 3'b000;
  assign _zz_46 = 3'b001;
  assign _zz_47 = 3'b001;
  assign _zz_48 = 3'b010;
  assign _zz_49 = 3'b001;
  assign _zz_50 = 3'b010;
  assign _zz_51 = 3'b010;
  assign _zz_52 = 3'b011;
  always @(*) begin
    LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id = LsuL1Plugin_logic_lsu_ctrl_wayId;
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_id = LsuL1Plugin_logic_lsu_ctrl_targetWay;
    end
  end

  assign LsuL1Plugin_logic_lsu_ctrl_doRefillPush = (LsuL1Plugin_logic_lsu_ctrl_doRefill || LsuL1Plugin_logic_lsu_ctrl_doUpgrade);
  always @(*) begin
    LsuL1Plugin_logic_refill_push_valid = LsuL1Plugin_logic_lsu_ctrl_doRefillPush;
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_refill_push_valid = 1'b0;
    end
  end

  assign LsuL1Plugin_logic_refill_push_payload_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign LsuL1Plugin_logic_refill_push_payload_unique = execute_ctrl4_down_LsuL1Plugin_logic_NEED_UNIQUE_lane0;
  assign LsuL1Plugin_logic_refill_push_payload_data = LsuL1Plugin_logic_lsu_ctrl_askRefill;
  always @(*) begin
    LsuL1Plugin_logic_refill_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_targetWay;
    if(LsuL1Plugin_logic_lsu_ctrl_askUpgrade) begin
      LsuL1Plugin_logic_refill_push_payload_way = LsuL1Plugin_logic_lsu_ctrl_wayId;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_refill_push_payload_victim = ((LsuL1Plugin_logic_lsu_ctrl_refillWayNeedWriteback && LsuL1Plugin_logic_lsu_ctrl_refillWayWasDirty) ? LsuL1Plugin_logic_writeback_free : 1'b0);
    if(LsuL1Plugin_logic_lsu_ctrl_askUpgrade) begin
      LsuL1Plugin_logic_refill_push_payload_victim = 1'b0;
    end
  end

  assign LsuL1Plugin_logic_refill_push_payload_dirty = execute_ctrl4_down_LsuL1_STORE_lane0;
  assign execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0 = (LsuL1Plugin_logic_lsu_ctrl_refillHazards | (((! execute_ctrl4_down_LsuL1_HAZARD_lane0) && (LsuL1Plugin_logic_lsu_ctrl_askRefill || LsuL1Plugin_logic_lsu_ctrl_askUpgrade)) ? (LsuL1Plugin_logic_refill_full ? 1'b1 : LsuL1Plugin_logic_refill_free) : 1'b0));
  assign execute_ctrl4_down_LsuL1_WAIT_WRITEBACK_lane0 = 1'b0;
  assign when_LsuL1Plugin_l915 = (execute_ctrl4_down_LsuL1_SEL_lane0 && (! execute_ctrl4_down_LsuL1_ABORD_lane0));
  assign _zz_53 = {LsuL1Plugin_logic_lsu_ctrl_askRefill,{LsuL1Plugin_logic_lsu_ctrl_doUpgrade,LsuL1Plugin_logic_lsu_ctrl_doFlush}};
  always @(*) begin
    LsuL1Plugin_logic_shared_write_valid = 1'b0;
    if(LsuL1Plugin_logic_lsu_ctrl_doFlush) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_doRefill) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(when_LsuL1Plugin_l1019) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
    if(LsuL1Plugin_logic_lsu_ctrl_preventSideEffects) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b0;
    end
    if(when_LsuL1Plugin_l1219) begin
      LsuL1Plugin_logic_shared_write_valid = 1'b1;
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_address = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0[11 : 6];
    if(when_LsuL1Plugin_l1219) begin
      LsuL1Plugin_logic_shared_write_payload_address = LsuL1Plugin_logic_initializer_counter[5:0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_data_plru_0 = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_0;
    if(when_LsuL1Plugin_l1219) begin
      LsuL1Plugin_logic_shared_write_payload_data_plru_0 = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0[0 : 0];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_data_plru_1 = LsuL1Plugin_logic_lsu_ctrl_plruLogic_core_io_update_state_1;
    if(when_LsuL1Plugin_l1219) begin
      LsuL1Plugin_logic_shared_write_payload_data_plru_1 = _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0[2 : 1];
    end
  end

  always @(*) begin
    LsuL1Plugin_logic_shared_write_payload_data_dirty = ((execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty | (LsuL1Plugin_logic_lsu_ctrl_doWrite ? execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 : 4'b0000)) & (~ ((LsuL1Plugin_logic_lsu_ctrl_doRefill ? _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty_1 : 4'b0000) | (LsuL1Plugin_logic_lsu_ctrl_doFlush ? LsuL1Plugin_logic_lsu_ctrl_needFlushOh : 4'b0000))));
    if(when_LsuL1Plugin_l1219) begin
      LsuL1Plugin_logic_shared_write_payload_data_dirty = _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty[6 : 3];
    end
  end

  assign _zz_54 = ({1'd0,1'b1} <<< execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0[2 : 2]);
  assign when_LsuL1Plugin_l929 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[0];
  assign when_LsuL1Plugin_l929_1 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[1];
  assign when_LsuL1Plugin_l929_2 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[2];
  assign when_LsuL1Plugin_l929_3 = execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0[3];
  assign execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0 = (|LsuL1Plugin_logic_lsu_ctrl_needFlushs);
  assign _zz_LsuL1Plugin_logic_waysWrite_tag_address = _zz__zz_LsuL1Plugin_logic_waysWrite_tag_address;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 = LsuL1Plugin_logic_lsu_ctrl_doWrite;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = execute_ctrl4_down_LsuL1_MASK_lane0;
  assign when_LsuL1Plugin_l1019 = ((execute_ctrl4_down_LsuL1_SEL_lane0 && (! execute_ctrl4_down_LsuL1_HAZARD_lane0)) && (! execute_ctrl4_down_LsuL1_MISS_lane0));
  always @(*) begin
    execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0 = execute_ctrl4_down_LsuL1Plugin_logic_MUXED_DATA_lane0;
    if(when_LsuL1Plugin_l1026) begin
      if(when_LsuL1Plugin_l1030) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[7 : 0] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[7 : 0];
      end
      if(when_LsuL1Plugin_l1030_1) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[15 : 8] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[15 : 8];
      end
      if(when_LsuL1Plugin_l1030_2) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[23 : 16] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[23 : 16];
      end
      if(when_LsuL1Plugin_l1030_3) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[31 : 24] = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[31 : 24];
      end
    end
    if(when_LsuL1Plugin_l1026_1) begin
      if(when_LsuL1Plugin_l1030_4) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[7 : 0] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[7 : 0];
      end
      if(when_LsuL1Plugin_l1030_5) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[15 : 8] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[15 : 8];
      end
      if(when_LsuL1Plugin_l1030_6) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[23 : 16] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[23 : 16];
      end
      if(when_LsuL1Plugin_l1030_7) begin
        execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0[31 : 24] = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0[31 : 24];
      end
    end
  end

  assign when_LsuL1Plugin_l1026 = execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[1];
  assign when_LsuL1Plugin_l1030 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[0];
  assign when_LsuL1Plugin_l1030_1 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[1];
  assign when_LsuL1Plugin_l1030_2 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[2];
  assign when_LsuL1Plugin_l1030_3 = execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[3];
  assign when_LsuL1Plugin_l1026_1 = execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0[0];
  assign when_LsuL1Plugin_l1030_4 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[0];
  assign when_LsuL1Plugin_l1030_5 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[1];
  assign when_LsuL1Plugin_l1030_6 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[2];
  assign when_LsuL1Plugin_l1030_7 = execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0[3];
  assign execute_ctrl4_down_LsuL1_READ_DATA_lane0 = execute_ctrl4_down_LsuL1Plugin_logic_BYPASSED_DATA_lane0;
  assign LsuL1Plugin_logic_initializer_done = LsuL1Plugin_logic_initializer_counter[6];
  assign when_LsuL1Plugin_l1219 = (! LsuL1Plugin_logic_initializer_done);
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty = 7'h0;
  assign _zz_LsuL1Plugin_logic_shared_write_payload_data_plru_0 = _zz_LsuL1Plugin_logic_shared_write_payload_data_dirty[2 : 0];
  assign LsuL1Plugin_logic_refill_read_reservation_win = (! 1'b0);
  assign LsuL1Plugin_logic_lsu_ctrl_wayWriteReservation_win = (! (|LsuL1Plugin_logic_refill_read_reservation_take));
  assign LsuL1Plugin_logic_refill_read_writeReservation_win = (! 1'b0);
  assign LsuL1Plugin_logic_lsu_ctrl_bankWriteReservation_win = (! (|LsuL1Plugin_logic_refill_read_writeReservation_take));
  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_address = 4'bxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_address = _zz_TrapPlugin_logic_harts_0_crsPorts_write_address;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_address = _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_crsPorts_write_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        TrapPlugin_logic_harts_0_crsPorts_write_data = TrapPlugin_logic_harts_0_trap_pending_pc;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        TrapPlugin_logic_harts_0_crsPorts_write_data = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval;
        if(TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg) begin
          TrapPlugin_logic_harts_0_crsPorts_write_data = TrapPlugin_logic_harts_0_trap_pending_pc;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_interrupt_valid = 1'b0;
    if(when_TrapPlugin_l201_1) begin
      if(when_TrapPlugin_l207) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l207_1) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l207_2) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
    end
    if(when_TrapPlugin_l201) begin
      if(when_TrapPlugin_l207_3) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l207_4) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l207_5) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l207_6) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l207_7) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
      if(when_TrapPlugin_l207_8) begin
        TrapPlugin_logic_harts_0_interrupt_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_interrupt_code = 4'bxxxx;
    if(when_TrapPlugin_l201_1) begin
      if(when_TrapPlugin_l207) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0001;
      end
      if(when_TrapPlugin_l207_1) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0101;
      end
      if(when_TrapPlugin_l207_2) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b1001;
      end
    end
    if(when_TrapPlugin_l201) begin
      if(when_TrapPlugin_l207_3) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0111;
      end
      if(when_TrapPlugin_l207_4) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0011;
      end
      if(when_TrapPlugin_l207_5) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b1011;
      end
      if(when_TrapPlugin_l207_6) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0001;
      end
      if(when_TrapPlugin_l207_7) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b0101;
      end
      if(when_TrapPlugin_l207_8) begin
        TrapPlugin_logic_harts_0_interrupt_code = 4'b1001;
      end
    end
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'bxx;
    if(when_TrapPlugin_l201_1) begin
      if(when_TrapPlugin_l207) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b01;
      end
      if(when_TrapPlugin_l207_1) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b01;
      end
      if(when_TrapPlugin_l207_2) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b01;
      end
    end
    if(when_TrapPlugin_l201) begin
      if(when_TrapPlugin_l207_3) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l207_4) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l207_5) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l207_6) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l207_7) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
      if(when_TrapPlugin_l207_8) begin
        TrapPlugin_logic_harts_0_interrupt_targetPrivilege = 2'b11;
      end
    end
  end

  assign when_TrapPlugin_l201 = (PrivilegedPlugin_logic_harts_0_m_status_mie || (! PrivilegedPlugin_logic_harts_0_withMachinePrivilege));
  assign when_TrapPlugin_l201_1 = ((PrivilegedPlugin_logic_harts_0_s_status_sie && (! PrivilegedPlugin_logic_harts_0_withMachinePrivilege)) || (! PrivilegedPlugin_logic_harts_0_withSupervisorPrivilege));
  assign when_TrapPlugin_l207 = ((_zz_when_TrapPlugin_l207_3 && (1'b1 && PrivilegedPlugin_logic_harts_0_m_ideleg_ss)) && (! 1'b0));
  assign when_TrapPlugin_l207_1 = ((_zz_when_TrapPlugin_l207_4 && (1'b1 && PrivilegedPlugin_logic_harts_0_m_ideleg_st)) && (! 1'b0));
  assign when_TrapPlugin_l207_2 = ((_zz_when_TrapPlugin_l207_5 && (1'b1 && PrivilegedPlugin_logic_harts_0_m_ideleg_se)) && (! 1'b0));
  assign when_TrapPlugin_l207_3 = ((_zz_when_TrapPlugin_l207 && 1'b1) && (! 1'b0));
  assign when_TrapPlugin_l207_4 = ((_zz_when_TrapPlugin_l207_1 && 1'b1) && (! 1'b0));
  assign when_TrapPlugin_l207_5 = ((_zz_when_TrapPlugin_l207_2 && 1'b1) && (! 1'b0));
  assign when_TrapPlugin_l207_6 = ((_zz_when_TrapPlugin_l207_3 && 1'b1) && (! (|PrivilegedPlugin_logic_harts_0_m_ideleg_ss)));
  assign when_TrapPlugin_l207_7 = ((_zz_when_TrapPlugin_l207_4 && 1'b1) && (! (|PrivilegedPlugin_logic_harts_0_m_ideleg_st)));
  assign when_TrapPlugin_l207_8 = ((_zz_when_TrapPlugin_l207_5 && 1'b1) && (! (|PrivilegedPlugin_logic_harts_0_m_ideleg_se)));
  assign TrapPlugin_logic_harts_0_interrupt_pendingInterrupt = (TrapPlugin_logic_harts_0_interrupt_validBuffer && PrivilegedPlugin_api_harts_0_allowInterrupts);
  assign when_TrapPlugin_l226 = (|{_zz_when_TrapPlugin_l207_5,{_zz_when_TrapPlugin_l207_4,{_zz_when_TrapPlugin_l207_3,{_zz_when_TrapPlugin_l207_2,{_zz_when_TrapPlugin_l207_1,_zz_when_TrapPlugin_l207}}}}});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid = (early0_EnvPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_valid = (FetchL1Plugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid = (LsuPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid = (early0_BranchPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1 = (CsrAccessPlugin_logic_trapPort_valid && 1'b1);
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid = (DecoderPlugin_logic_laneLogic_0_trapPort_valid && 1'b1);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_exception = LsuPlugin_logic_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_tval = LsuPlugin_logic_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_code = LsuPlugin_logic_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg = LsuPlugin_logic_trapPort_payload_arg;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_exception = early0_BranchPlugin_logic_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_tval = early0_BranchPlugin_logic_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_code = early0_BranchPlugin_logic_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg = early0_BranchPlugin_logic_trapPort_payload_arg;
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception = {(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1 && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid && 1'b0)))),(_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid && (&(! (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1 && 1'b0))))};
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1 = ((_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception[0] ? {early0_EnvPlugin_logic_trapPort_payload_arg,{early0_EnvPlugin_logic_trapPort_payload_code,{early0_EnvPlugin_logic_trapPort_payload_tval,early0_EnvPlugin_logic_trapPort_payload_exception}}} : 40'h0) | (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception[1] ? {CsrAccessPlugin_logic_trapPort_payload_arg,{CsrAccessPlugin_logic_trapPort_payload_code,{CsrAccessPlugin_logic_trapPort_payload_tval,CsrAccessPlugin_logic_trapPort_payload_exception}}} : 40'h0));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[32 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[36 : 33];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_exception_1[39 : 37];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_exception = DecoderPlugin_logic_laneLogic_0_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_tval = DecoderPlugin_logic_laneLogic_0_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_code = DecoderPlugin_logic_laneLogic_0_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg = DecoderPlugin_logic_laneLogic_0_trapPort_payload_arg;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_valid = (|_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_valid);
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_exception = FetchL1Plugin_logic_trapPort_payload_exception;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_tval = FetchL1Plugin_logic_trapPort_payload_tval;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_code = FetchL1Plugin_logic_trapPort_payload_code;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_arg = FetchL1Plugin_logic_trapPort_payload_arg;
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh = {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_valid,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid,TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid}}}};
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[0];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[1];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[2];
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4 = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[3];
  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_5[0] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1 && (! 1'b0));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_5[1] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2 && (! _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_5[2] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3 && (! (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1})));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_5[3] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4 && (! (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1}})));
    _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_5[4] = (_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[4] && (! (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_4,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_3,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_2,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_1}}})));
  end

  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_oh = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_oh_5;
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid = (|{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_valid,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid_1,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_valid,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_valid,{_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_valid,_zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_valid}}}}});
  assign _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = ((((TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[0] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_0_payload_arg,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception} : 40'h0) | (TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[1] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_1_payload_arg,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_1} : 40'h0)) | ((TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[2] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_2_payload_arg,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_2} : 40'h0) | (TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[3] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_3_payload_arg,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_3} : 40'h0))) | (TrapPlugin_logic_harts_0_trap_pending_arbiter_oh[4] ? {TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_arg,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_code,{TrapPlugin_logic_harts_0_trap_pending_arbiter_ports_4_payload_tval,_zz__zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception_4}}} : 40'h0));
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[0];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[32 : 1];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[36 : 33];
  assign TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg = _zz_TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception[39 : 37];
  assign TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege = PrivilegedPlugin_logic_harts_0_m_status_mpp;
    case(TrapPlugin_logic_harts_0_trap_pending_xret_sourcePrivilege)
      2'b01 : begin
        TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege = {1'b0,PrivilegedPlugin_logic_harts_0_s_status_spp};
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b11;
    case(TrapPlugin_logic_harts_0_trap_exception_code)
      4'b0000 : begin
        if(when_TrapPlugin_l263) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b0011 : begin
        if(when_TrapPlugin_l263_1) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1000 : begin
        if(when_TrapPlugin_l263_2) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1001 : begin
        if(when_TrapPlugin_l263_3) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1100 : begin
        if(when_TrapPlugin_l263_4) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1101 : begin
        if(when_TrapPlugin_l263_5) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      4'b1111 : begin
        if(when_TrapPlugin_l263_6) begin
          TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped = 2'b01;
        end
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_exception_code = TrapPlugin_logic_harts_0_trap_pending_state_code;
  assign when_TrapPlugin_l263 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_iam) && (! 1'b0));
  assign when_TrapPlugin_l263_1 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_bp) && (! 1'b0));
  assign when_TrapPlugin_l263_2 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_eu) && (! 1'b0));
  assign when_TrapPlugin_l263_3 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_es) && (! 1'b0));
  assign when_TrapPlugin_l263_4 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_ipf) && (! 1'b0));
  assign when_TrapPlugin_l263_5 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_lpf) && (! 1'b0));
  assign when_TrapPlugin_l263_6 = ((1'b1 && PrivilegedPlugin_logic_harts_0_m_edeleg_spf) && (! 1'b0));
  assign TrapPlugin_logic_harts_0_trap_exception_targetPrivilege = ((PrivilegedPlugin_logic_harts_0_privilege < TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped) ? TrapPlugin_logic_harts_0_trap_exception_exceptionTargetPrivilegeUncapped : PrivilegedPlugin_logic_harts_0_privilege);
  assign PrivilegedPlugin_logic_harts_0_commitMask = (((execute_ctrl5_down_LANE_SEL_lane0 && execute_ctrl5_down_isReady) && (! execute_lane0_ctrls_5_downIsCancel)) && execute_ctrl5_down_COMMIT_lane0);
  assign TrapPlugin_logic_harts_0_trap_trigger_oh = (((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_TRAP_lane0);
  assign TrapPlugin_logic_harts_0_trap_trigger_valid = (|TrapPlugin_logic_harts_0_trap_trigger_oh);
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_trap = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_trap = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_interrupt = 1'bx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_interrupt = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_whitebox_code = 4'bxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_whitebox_code = TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_historyPort_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
        TrapPlugin_logic_harts_0_trap_historyPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_historyPort_payload_history = TrapPlugin_logic_harts_0_trap_pending_history;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        TrapPlugin_logic_harts_0_trap_pcPort_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_pcPort_payload_fault = 1'b0;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_pending_pc;
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_readed;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_readed;
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        TrapPlugin_logic_harts_0_trap_pcPort_payload_pc = TrapPlugin_logic_harts_0_trap_fsm_jumpTarget;
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_wantExit = 1'b0;
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_wantStart = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
        TrapPlugin_logic_harts_0_trap_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_wantKill = 1'b0;
  assign TrapPlugin_logic_harts_0_trap_fsm_inflightTrap = (|{execute_lane0_logic_trapPending[0],{DispatchPlugin_logic_trapPendings[0],decode_logic_trapPending[0]}});
  assign TrapPlugin_logic_harts_0_trap_fsm_holdPort = (TrapPlugin_logic_harts_0_trap_fsm_inflightTrap || (! (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RUNNING)));
  assign TrapPlugin_api_harts_0_fsmBusy = (! (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RUNNING));
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_wfi = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
              TrapPlugin_logic_harts_0_trap_fsm_wfi = 1'b1;
            end
            4'b0110 : begin
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
        if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt = 1'b1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt = ((TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0000) && TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege = (TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt ? TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege : TrapPlugin_logic_harts_0_trap_exception_targetPrivilege);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_tval = ((! TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt) ? TrapPlugin_logic_harts_0_trap_pending_state_tval : 32'h0);
  assign TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code = (TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt ? TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code : TrapPlugin_logic_harts_0_trap_pending_state_code);
  assign TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0 = (! TrapPlugin_logic_initHold);
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
            end
            4'b0111 : begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_valid = 1'b1;
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_address = TrapPlugin_logic_harts_0_trap_pending_state_tval;
  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_payload_storageId = TrapPlugin_logic_harts_0_trap_pending_state_arg[2 : 2];
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid = 1'b0;
    if(when_TrapPlugin_l355) begin
      TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid = 1'b1;
    end
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
        if(!when_TrapPlugin_l409) begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
            end
            4'b0001 : begin
            end
            4'b0010 : begin
            end
            4'b0100 : begin
            end
            4'b0101 : begin
            end
            4'b1000 : begin
            end
            4'b0110 : begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid = 1'b1;
            end
            4'b0111 : begin
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_fire = (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_valid && TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready);
  assign when_TrapPlugin_l355 = (! TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated);
  assign TrapPlugin_logic_harts_0_trap_fsm_jumpOffset = ((|{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b1000),{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0110),{(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0010),(TrapPlugin_logic_harts_0_trap_pending_state_code == 4'b0101)}}}) ? TrapPlugin_logic_harts_0_trap_pending_slices : 1'b0);
  always @(*) begin
    TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
        TrapPlugin_logic_fetchL1Invalidate_0_cmd_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid = 1'b0;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
        TrapPlugin_logic_lsuL1Invalidate_0_cmd_valid = 1'b1;
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak = 1'b0;
  assign when_TrapPlugin_l556 = (TrapPlugin_logic_harts_0_crsPorts_read_valid && TrapPlugin_logic_harts_0_crsPorts_read_ready);
  assign TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  always @(*) begin
    LsuPlugin_logic_flusher_arbiter_io_output_ready = 1'b0;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_CMD : begin
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
        if(when_LsuPlugin_l371) begin
          LsuPlugin_logic_flusher_arbiter_io_output_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign PrivilegedPlugin_api_lsuTriggerBus_load = execute_ctrl3_down_LsuL1_LOAD_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_store = execute_ctrl3_down_LsuL1_STORE_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_virtual = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
  assign PrivilegedPlugin_api_lsuTriggerBus_size = execute_ctrl3_down_LsuL1_SIZE_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0 = 1'b0;
  assign execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0 = (execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0 || execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0);
  assign LsuPlugin_logic_onAddress0_ls_prefetchOp = execute_ctrl2_down_Decode_UOP_lane0[24 : 20];
  assign LsuPlugin_logic_onAddress0_ls_port_valid = (execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_AguPlugin_SEL_lane0);
  assign LsuPlugin_logic_onAddress0_ls_port_payload_address = execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_size = execute_ctrl2_down_AguPlugin_SIZE_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_load = execute_ctrl2_down_AguPlugin_LOAD_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_store = execute_ctrl2_down_AguPlugin_STORE_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_atomic = execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_clean = 1'b0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_invalidate = 1'b0;
  assign LsuPlugin_logic_onAddress0_ls_port_payload_op = LsuL1CmdOpcode_LSU;
  assign LsuPlugin_logic_onAddress0_ls_port_fire = (LsuPlugin_logic_onAddress0_ls_port_valid && LsuPlugin_logic_onAddress0_ls_port_ready);
  assign LsuPlugin_logic_onAddress0_ls_port_payload_storeId = LsuPlugin_logic_onAddress0_ls_storeId;
  assign when_LsuPlugin_l259 = (|(LsuPlugin_logic_onAddress0_access_waiter_refill & (~ LsuL1_REFILL_BUSY)));
  assign LsuPlugin_logic_onAddress0_access_sbWaiter = 1'b0;
  assign _zz_MmuPlugin_logic_accessBus_cmd_ready = (! (LsuPlugin_logic_onAddress0_access_waiter_valid || LsuPlugin_logic_onAddress0_access_sbWaiter));
  assign MmuPlugin_logic_accessBus_cmd_haltWhen_valid = (MmuPlugin_logic_accessBus_cmd_valid && _zz_MmuPlugin_logic_accessBus_cmd_ready);
  assign MmuPlugin_logic_accessBus_cmd_ready = (MmuPlugin_logic_accessBus_cmd_haltWhen_ready && _zz_MmuPlugin_logic_accessBus_cmd_ready);
  assign MmuPlugin_logic_accessBus_cmd_haltWhen_payload_address = MmuPlugin_logic_accessBus_cmd_payload_address;
  assign MmuPlugin_logic_accessBus_cmd_haltWhen_payload_size = MmuPlugin_logic_accessBus_cmd_payload_size;
  assign LsuPlugin_logic_onAddress0_access_port_valid = MmuPlugin_logic_accessBus_cmd_haltWhen_valid;
  assign MmuPlugin_logic_accessBus_cmd_haltWhen_ready = LsuPlugin_logic_onAddress0_access_port_ready;
  assign LsuPlugin_logic_onAddress0_access_port_payload_address = MmuPlugin_logic_accessBus_cmd_payload_address;
  assign LsuPlugin_logic_onAddress0_access_port_payload_size = MmuPlugin_logic_accessBus_cmd_payload_size;
  assign LsuPlugin_logic_onAddress0_access_port_payload_load = 1'b1;
  assign LsuPlugin_logic_onAddress0_access_port_payload_store = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_atomic = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_clean = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_invalidate = 1'b0;
  assign LsuPlugin_logic_onAddress0_access_port_payload_op = LsuL1CmdOpcode_ACCESS_1;
  assign LsuPlugin_logic_onAddress0_access_port_payload_storeId = 12'h0;
  assign LsuPlugin_logic_onAddress0_flush_port_valid = ((LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_CMD) && (! LsuPlugin_logic_flusher_cmdCounter[6]));
  assign LsuPlugin_logic_onAddress0_flush_port_payload_address = {19'd0, _zz_LsuPlugin_logic_onAddress0_flush_port_payload_address};
  assign LsuPlugin_logic_onAddress0_flush_port_payload_size = 2'b00;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_load = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_store = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_atomic = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_clean = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_invalidate = 1'b0;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_op = LsuL1CmdOpcode_FLUSH;
  assign LsuPlugin_logic_onAddress0_flush_port_payload_storeId = 12'h0;
  assign LsuPlugin_logic_onAddress0_flush_port_fire = (LsuPlugin_logic_onAddress0_flush_port_valid && LsuPlugin_logic_onAddress0_flush_port_ready);
  assign LsuPlugin_logic_onAddress0_ls_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_0_ready;
  assign LsuPlugin_logic_onAddress0_access_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_1_ready;
  assign LsuPlugin_logic_onAddress0_flush_port_ready = LsuPlugin_logic_onAddress0_arbiter_io_inputs_2_ready;
  assign LsuPlugin_logic_onAddress0_arbiter_io_output_ready = (! execute_freeze_valid);
  assign execute_ctrl2_down_LsuL1_SEL_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_valid;
  assign execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address;
  always @(*) begin
    _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 4'bxxxx;
    case(LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size)
      2'b00 : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 4'b0001;
      end
      2'b01 : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 4'b0011;
      end
      2'b10 : begin
        _zz_execute_ctrl2_down_LsuL1_MASK_lane0 = 4'b1111;
      end
      default : begin
      end
    endcase
  end

  assign execute_ctrl2_down_LsuL1_MASK_lane0 = (_zz_execute_ctrl2_down_LsuL1_MASK_lane0 <<< LsuPlugin_logic_onAddress0_arbiter_io_output_payload_address[1 : 0]);
  assign execute_ctrl2_down_LsuL1_SIZE_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_size;
  assign execute_ctrl2_down_LsuL1_LOAD_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_load;
  assign execute_ctrl2_down_LsuL1_ATOMIC_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_atomic;
  assign execute_ctrl2_down_LsuL1_STORE_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_store;
  assign execute_ctrl2_down_LsuL1_CLEAN_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_clean;
  assign execute_ctrl2_down_LsuL1_INVALID_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_invalidate;
  assign execute_ctrl2_down_LsuL1_PREFETCH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_PREFETCH);
  assign execute_ctrl2_down_LsuL1_FLUSH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_FLUSH);
  assign execute_ctrl2_down_Decode_STORE_ID_lane0 = LsuPlugin_logic_onAddress0_arbiter_io_output_payload_storeId;
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_ACCESS_1);
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_WB_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_STORE_BUFFER);
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_LSU);
  assign execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = (LsuPlugin_logic_onAddress0_arbiter_io_output_payload_op == LsuL1CmdOpcode_PREFETCH);
  assign execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0 = execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign when_LsuPlugin_l546 = (execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 && (! execute_ctrl3_up_LANE_SEL_lane0));
  assign when_LsuPlugin_l546_1 = (execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (! execute_ctrl4_up_LANE_SEL_lane0));
  assign execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 = (|{((execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b10) && (execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[1 : 0] != 2'b00)),((execute_ctrl3_down_LsuL1_SIZE_lane0 == 2'b01) && (execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[0 : 0] != 1'b0))});
  assign execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0 = (((execute_ctrl3_down_AguPlugin_SEL_lane0 && execute_ctrl3_down_LsuL1_ATOMIC_lane0) && execute_ctrl3_down_LsuL1_STORE_lane0) && execute_ctrl3_down_LsuL1_LOAD_lane0);
  assign LsuPlugin_logic_onPma_cached_cmd_address = execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign LsuPlugin_logic_onPma_cached_cmd_op[0] = execute_ctrl3_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_address = execute_ctrl3_down_MMU_TRANSLATED_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_size = execute_ctrl3_down_LsuL1_SIZE_lane0;
  assign LsuPlugin_logic_onPma_io_cmd_op[0] = execute_ctrl3_down_LsuL1_STORE_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault = LsuPlugin_logic_onPma_cached_rsp_fault;
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io = LsuPlugin_logic_onPma_cached_rsp_io;
  always @(*) begin
    execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = LsuPlugin_logic_onPma_io_rsp_fault;
    if(when_LsuPlugin_l569) begin
      execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = 1'b1;
    end
  end

  assign execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io = LsuPlugin_logic_onPma_io_rsp_io;
  assign when_LsuPlugin_l569 = (execute_ctrl3_down_LsuL1_ATOMIC_lane0 || execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0);
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0 = (((execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault && (! execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault)) && (! execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0)) && (! execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0));
  assign LsuPlugin_logic_onPma_addressExtension = (MmuPlugin_api_lsuTranslationEnable ? _zz_LsuPlugin_logic_onPma_addressExtension[31] : 1'b0);
  assign execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = (execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 && 1'b0);
  assign execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 = (execute_ctrl3_down_MMU_PAGE_FAULT_lane0 || (execute_ctrl3_down_AguPlugin_STORE_lane0 ? (! execute_ctrl3_down_MMU_ALLOW_WRITE_lane0) : (! execute_ctrl3_down_MMU_ALLOW_READ_lane0)));
  assign execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0 = ((((execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 || execute_ctrl3_down_MMU_ACCESS_FAULT_lane0) || execute_ctrl3_down_MMU_REFILL_lane0) || execute_ctrl3_down_MMU_HAZARD_lane0) || execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0);
  always @(*) begin
    LsuPlugin_logic_onCtrl_lsuTrap = 1'b0;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b1;
    end
    if(when_LsuPlugin_l833) begin
      LsuPlugin_logic_onCtrl_lsuTrap = 1'b0;
    end
  end

  always @(*) begin
    LsuPlugin_logic_onCtrl_writeData = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    LsuPlugin_logic_onCtrl_writeData[31 : 0] = execute_ctrl4_up_integer_RS2_lane0;
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0) begin
      LsuPlugin_logic_onCtrl_writeData[31 : 0] = LsuPlugin_logic_onCtrl_rva_aluBuffer;
    end
  end

  assign when_LsuPlugin_l597 = (((((! LsuPlugin_logic_onCtrl_lsuTrap) && (! execute_lane0_ctrls_4_upIsCancel)) && execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0) && (! execute_ctrl4_down_LsuL1_CLEAN_lane0)) && (! execute_ctrl4_down_LsuL1_INVALID_lane0));
  assign LsuPlugin_logic_onCtrl_io_doIt = ((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_LsuL1_SEL_lane0) && execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0);
  assign LsuPlugin_logic_bus_cmd_fire = (LsuPlugin_logic_bus_cmd_valid && LsuPlugin_logic_bus_cmd_ready);
  assign when_LsuPlugin_l601 = (! execute_freeze_valid);
  assign LsuPlugin_logic_bus_cmd_valid = (((LsuPlugin_logic_onCtrl_io_doItReg && (! LsuPlugin_logic_onCtrl_io_cmdSent)) && LsuPlugin_logic_onCtrl_io_allowIt) && (! LsuPlugin_logic_onCtrl_io_tooEarly));
  assign LsuPlugin_logic_bus_cmd_payload_write = execute_ctrl4_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_data = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_size = execute_ctrl4_down_LsuL1_SIZE_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_mask = execute_ctrl4_down_LsuL1_MASK_lane0;
  assign LsuPlugin_logic_bus_cmd_payload_io = 1'b1;
  assign LsuPlugin_logic_bus_cmd_payload_fromHart = 1'b1;
  assign LsuPlugin_logic_bus_cmd_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign LsuPlugin_logic_bus_rsp_toStream_valid = LsuPlugin_logic_bus_rsp_valid;
  assign LsuPlugin_logic_bus_rsp_toStream_payload_error = LsuPlugin_logic_bus_rsp_payload_error;
  assign LsuPlugin_logic_bus_rsp_toStream_payload_data = LsuPlugin_logic_bus_rsp_payload_data;
  assign LsuPlugin_logic_onCtrl_io_rsp_fire = (LsuPlugin_logic_onCtrl_io_rsp_valid && LsuPlugin_logic_onCtrl_io_rsp_ready);
  assign LsuPlugin_logic_bus_rsp_toStream_ready = (! LsuPlugin_logic_bus_rsp_toStream_rValid);
  assign LsuPlugin_logic_onCtrl_io_rsp_valid = LsuPlugin_logic_bus_rsp_toStream_rValid;
  assign LsuPlugin_logic_onCtrl_io_rsp_payload_error = LsuPlugin_logic_bus_rsp_toStream_rData_error;
  assign LsuPlugin_logic_onCtrl_io_rsp_payload_data = LsuPlugin_logic_bus_rsp_toStream_rData_data;
  assign LsuPlugin_logic_onCtrl_io_rsp_ready = (! execute_freeze_valid);
  assign LsuPlugin_logic_onCtrl_io_freezeIt = (LsuPlugin_logic_onCtrl_io_doIt && (LsuPlugin_logic_onCtrl_io_tooEarly || ((! LsuPlugin_logic_onCtrl_io_rsp_valid) && LsuPlugin_logic_onCtrl_io_allowIt)));
  assign LsuPlugin_logic_onCtrl_loadData_input = (LsuPlugin_logic_onCtrl_io_cmdSent ? LsuPlugin_logic_onCtrl_io_rsp_payload_data : execute_ctrl4_down_LsuL1_READ_DATA_lane0);
  assign LsuPlugin_logic_onCtrl_loadData_splitted_0 = LsuPlugin_logic_onCtrl_loadData_input[7 : 0];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_1 = LsuPlugin_logic_onCtrl_loadData_input[15 : 8];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_2 = LsuPlugin_logic_onCtrl_loadData_input[23 : 16];
  assign LsuPlugin_logic_onCtrl_loadData_splitted_3 = LsuPlugin_logic_onCtrl_loadData_input[31 : 24];
  always @(*) begin
    LsuPlugin_logic_onCtrl_loadData_shifted[7 : 0] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted;
    LsuPlugin_logic_onCtrl_loadData_shifted[15 : 8] = _zz_LsuPlugin_logic_onCtrl_loadData_shifted_2;
    LsuPlugin_logic_onCtrl_loadData_shifted[23 : 16] = LsuPlugin_logic_onCtrl_loadData_splitted_2;
    LsuPlugin_logic_onCtrl_loadData_shifted[31 : 24] = LsuPlugin_logic_onCtrl_loadData_splitted_3;
  end

  assign execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0 = LsuPlugin_logic_onCtrl_loadData_shifted;
  assign LsuPlugin_logic_onCtrl_storeData_mapping_0_1 = {4{LsuPlugin_logic_onCtrl_writeData[7 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_1_1 = {2{LsuPlugin_logic_onCtrl_writeData[15 : 0]}};
  assign LsuPlugin_logic_onCtrl_storeData_mapping_2_1 = {1{LsuPlugin_logic_onCtrl_writeData[31 : 0]}};
  always @(*) begin
    _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(execute_ctrl4_down_LsuL1_SIZE_lane0)
      2'b00 : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_0_1;
      end
      2'b01 : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_1_1;
      end
      2'b10 : begin
        _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = LsuPlugin_logic_onCtrl_storeData_mapping_2_1;
      end
      default : begin
      end
    endcase
  end

  assign execute_ctrl4_down_LsuL1_WRITE_DATA_lane0 = _zz_execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0 = LsuPlugin_logic_onCtrl_scMiss;
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_compare = execute_ctrl4_down_Decode_UOP_lane0[31 : 29];
  assign _zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf = execute_ctrl4_down_Decode_UOP_lane0[27];
  assign LsuPlugin_logic_onCtrl_rva_alu_compare = _zz_LsuPlugin_logic_onCtrl_rva_alu_compare[2];
  assign LsuPlugin_logic_onCtrl_rva_alu_unsigned = _zz_LsuPlugin_logic_onCtrl_rva_alu_compare[1];
  assign LsuPlugin_logic_onCtrl_rva_alu_addSub = _zz_LsuPlugin_logic_onCtrl_rva_alu_addSub;
  assign LsuPlugin_logic_onCtrl_rva_alu_less = ((execute_ctrl4_down_integer_RS2_lane0[31] == LsuPlugin_logic_onCtrl_rva_srcBuffer[31]) ? LsuPlugin_logic_onCtrl_rva_alu_addSub[31] : (LsuPlugin_logic_onCtrl_rva_alu_unsigned ? LsuPlugin_logic_onCtrl_rva_srcBuffer[31] : execute_ctrl4_down_integer_RS2_lane0[31]));
  assign LsuPlugin_logic_onCtrl_rva_alu_selectRf = (_zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf ? 1'b1 : (_zz_LsuPlugin_logic_onCtrl_rva_alu_compare[0] ^ LsuPlugin_logic_onCtrl_rva_alu_less));
  assign switch_Misc_l242_1 = (_zz_LsuPlugin_logic_onCtrl_rva_alu_compare | {_zz_LsuPlugin_logic_onCtrl_rva_alu_selectRf,2'b00});
  always @(*) begin
    case(switch_Misc_l242_1)
      3'b000 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = LsuPlugin_logic_onCtrl_rva_alu_addSub;
      end
      3'b001 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (execute_ctrl4_down_integer_RS2_lane0 ^ LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      3'b010 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (execute_ctrl4_down_integer_RS2_lane0 | LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      3'b011 : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (execute_ctrl4_down_integer_RS2_lane0 & LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
      default : begin
        LsuPlugin_logic_onCtrl_rva_alu_raw = (LsuPlugin_logic_onCtrl_rva_alu_selectRf ? execute_ctrl4_down_integer_RS2_lane0 : LsuPlugin_logic_onCtrl_rva_srcBuffer);
      end
    endcase
  end

  assign LsuPlugin_logic_onCtrl_rva_alu_result = LsuPlugin_logic_onCtrl_rva_alu_raw;
  assign LsuPlugin_logic_onCtrl_rva_delay_0 = _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
  assign LsuPlugin_logic_onCtrl_rva_delay_1 = _zz_LsuPlugin_logic_onCtrl_rva_delay_1;
  assign LsuPlugin_logic_onCtrl_rva_freezeIt = ((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0) && (|{LsuPlugin_logic_onCtrl_rva_delay_1,LsuPlugin_logic_onCtrl_rva_delay_0}));
  always @(*) begin
    LsuPlugin_logic_onCtrl_rva_lrsc_capture = 1'b0;
    if(when_LsuPlugin_l685) begin
      if(!execute_ctrl4_down_LsuL1_STORE_lane0) begin
        if(execute_ctrl4_down_LsuL1_ATOMIC_lane0) begin
          LsuPlugin_logic_onCtrl_rva_lrsc_capture = 1'b1;
        end
      end
    end
  end

  assign when_LsuPlugin_l685 = ((((((! execute_freeze_valid) && execute_ctrl4_up_LANE_SEL_lane0) && execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0) && execute_ctrl4_down_LsuL1_SEL_lane0) && (! LsuPlugin_logic_onCtrl_lsuTrap)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0));
  assign LsuPlugin_logic_onCtrl_scMiss = (! LsuPlugin_logic_onCtrl_rva_lrsc_reserved);
  assign LsuL1_lockPort_valid = LsuPlugin_logic_onCtrl_rva_lrsc_reserved;
  assign LsuL1_lockPort_address = LsuPlugin_logic_onCtrl_rva_lrsc_address;
  assign when_LsuPlugin_l697 = (LsuPlugin_logic_onCtrl_rva_lrsc_age[5] || LsuPlugin_logic_onCtrl_io_cmdSent);
  always @(*) begin
    LsuPlugin_logic_flushPort_valid = 1'b0;
    if(when_LsuPlugin_l861) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        LsuPlugin_logic_flushPort_valid = 1'b1;
      end
    end
  end

  assign LsuPlugin_logic_flushPort_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign LsuPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    LsuPlugin_logic_trapPort_valid = 1'b0;
    if(when_LsuPlugin_l861) begin
      if(LsuPlugin_logic_onCtrl_lsuTrap) begin
        LsuPlugin_logic_trapPort_valid = 1'b1;
      end
    end
  end

  assign LsuPlugin_logic_trapPort_payload_tval = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  always @(*) begin
    LsuPlugin_logic_trapPort_payload_exception = 1'bx;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b1;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_trapPort_payload_exception = 1'b0;
    end
  end

  always @(*) begin
    LsuPlugin_logic_trapPort_payload_code = 4'bxxxx;
    if(LsuPlugin_logic_onCtrl_traps_accessFault) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(LsuPlugin_logic_onCtrl_traps_l1Failed) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b1101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(execute_ctrl4_down_MMU_ACCESS_FAULT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
    end
    if(execute_ctrl4_down_MMU_REFILL_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0111;
    end
    if(execute_ctrl4_down_MMU_HAZARD_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0100;
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0101;
      if(execute_ctrl4_down_AguPlugin_STORE_lane0) begin
        LsuPlugin_logic_trapPort_payload_code[1] = 1'b1;
      end
      if(when_LsuPlugin_l806) begin
        LsuPlugin_logic_trapPort_payload_code[3] = 1'b1;
      end
    end
    if(execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = {1'd0, _zz_LsuPlugin_logic_trapPort_payload_code};
    end
    if(execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0) begin
      LsuPlugin_logic_trapPort_payload_code = 4'b0011;
    end
  end

  always @(*) begin
    LsuPlugin_logic_trapPort_payload_arg = 3'b000;
    LsuPlugin_logic_trapPort_payload_arg[1 : 0] = (execute_ctrl4_down_LsuL1_STORE_lane0 ? 2'b01 : 2'b00);
    LsuPlugin_logic_trapPort_payload_arg[2 : 2] = 1'b1;
  end

  assign LsuPlugin_logic_onCtrl_traps_accessFault = ((execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault ? (LsuPlugin_logic_onCtrl_io_rsp_valid && LsuPlugin_logic_onCtrl_io_rsp_payload_error) : execute_ctrl4_down_LsuL1_FAULT_lane0) || execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0);
  assign LsuPlugin_logic_onCtrl_traps_l1Failed = ((! execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault) && (execute_ctrl4_down_LsuL1_HAZARD_lane0 || ((execute_ctrl4_down_LsuL1_MISS_lane0 || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0) && (execute_ctrl4_down_LsuL1_LOAD_lane0 || execute_ctrl4_down_LsuL1_STORE_lane0))));
  assign LsuPlugin_logic_onCtrl_traps_pmaFault = (execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault && execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault);
  assign when_LsuPlugin_l806 = (! execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0);
  assign when_LsuPlugin_l833 = (execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0 || execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0);
  assign when_LsuPlugin_l861 = (execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_AguPlugin_SEL_lane0);
  assign LsuPlugin_logic_onCtrl_mmuNeeded = (execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 || execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0);
  assign execute_ctrl4_down_LsuL1_ABORD_lane0 = (|{(LsuPlugin_logic_onCtrl_mmuNeeded && execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0),{(execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (((! execute_ctrl4_up_LANE_SEL_lane0) || execute_lane0_ctrls_4_upIsCancel) || execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0)),{((! execute_ctrl4_down_LsuL1_FLUSH_lane0) && execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault),{execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0,execute_ctrl4_down_LsuL1_HAZARD_lane0}}}});
  assign execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0 = (|{((execute_ctrl4_down_LsuL1_ATOMIC_lane0 && (! execute_ctrl4_down_LsuL1_LOAD_lane0)) && LsuPlugin_logic_onCtrl_scMiss),{execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0,{(execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 && (execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0 || execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0)),{execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0,{execute_ctrl4_down_LsuL1_FAULT_lane0,(execute_ctrl4_down_LsuL1_MISS_lane0 || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0)}}}}});
  assign when_LsuPlugin_l901 = ((execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuL1_FLUSH_lane0) && ((execute_ctrl4_down_LsuL1_FLUSH_HIT_lane0 || execute_ctrl4_down_LsuL1_HAZARD_lane0) || execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0));
  assign MmuPlugin_logic_accessBus_rsp_valid = ((execute_ctrl4_down_LsuL1_SEL_lane0 && execute_ctrl4_down_LsuPlugin_logic_FROM_ACCESS_lane0) && (! execute_freeze_valid));
  assign MmuPlugin_logic_accessBus_rsp_payload_data = execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
  always @(*) begin
    MmuPlugin_logic_accessBus_rsp_payload_error = (execute_ctrl4_down_LsuL1_FAULT_lane0 || execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0);
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      MmuPlugin_logic_accessBus_rsp_payload_error = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_logic_accessBus_rsp_payload_redo = LsuPlugin_logic_onCtrl_traps_l1Failed;
    if(LsuPlugin_logic_onCtrl_traps_pmaFault) begin
      MmuPlugin_logic_accessBus_rsp_payload_redo = 1'b0;
    end
  end

  assign MmuPlugin_logic_accessBus_rsp_payload_waitAny = 1'b0;
  assign when_LsuPlugin_l938 = (MmuPlugin_logic_accessBus_rsp_valid && MmuPlugin_logic_accessBus_rsp_payload_redo);
  assign when_LsuPlugin_l263 = (|execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0);
  assign when_LsuPlugin_l259_1 = (|(LsuPlugin_logic_onCtrl_hartRegulation_refill & (~ LsuL1_REFILL_BUSY)));
  assign when_LsuPlugin_l945 = ((((((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_down_AguPlugin_SEL_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0)) && 1'b1) && ((execute_ctrl4_down_LsuL1_HAZARD_lane0 || execute_ctrl4_down_LsuL1_MISS_lane0) || execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0));
  assign when_LsuPlugin_l263_1 = (|execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0);
  assign LsuPlugin_logic_commitProbe_valid = (((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && (execute_ctrl4_down_AguPlugin_SEL_lane0 ? execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 : (execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0 && execute_ctrl4_down_LsuL1_HAZARD_lane0)));
  assign LsuPlugin_logic_commitProbe_payload_address = execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0;
  assign LsuPlugin_logic_commitProbe_payload_load = execute_ctrl4_down_LsuL1_LOAD_lane0;
  assign LsuPlugin_logic_commitProbe_payload_store = execute_ctrl4_down_LsuL1_STORE_lane0;
  assign LsuPlugin_logic_commitProbe_payload_trap = LsuPlugin_logic_onCtrl_lsuTrap;
  assign LsuPlugin_logic_commitProbe_payload_miss = ((execute_ctrl4_down_LsuL1_MISS_lane0 && (! execute_ctrl4_down_LsuL1_HAZARD_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0));
  assign LsuPlugin_logic_commitProbe_payload_io = execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0;
  assign LsuPlugin_logic_commitProbe_payload_prefetchFailed = execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign LsuPlugin_logic_commitProbe_payload_pc = execute_ctrl4_down_PC_lane0;
  assign LsuPlugin_logic_iwb_valid = (execute_ctrl4_down_AguPlugin_SEL_lane0 && (! execute_ctrl4_down_AguPlugin_FLOAT_lane0));
  always @(*) begin
    LsuPlugin_logic_iwb_payload = execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
    if(when_LsuPlugin_l968) begin
      LsuPlugin_logic_iwb_payload[0] = execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
      LsuPlugin_logic_iwb_payload[7 : 1] = 7'h0;
    end
  end

  assign when_LsuPlugin_l968 = (execute_ctrl4_down_LsuL1_ATOMIC_lane0 && (! execute_ctrl4_down_LsuL1_LOAD_lane0));
  assign LsuPlugin_logic_onWb_storeFire = ((((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && execute_ctrl4_down_LsuL1_STORE_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0));
  assign LsuPlugin_logic_onWb_storeBroadcast = (((((((execute_ctrl4_down_isReady && execute_ctrl4_down_LsuL1_SEL_lane0) && execute_ctrl4_down_LsuL1_STORE_lane0) && (! execute_ctrl4_down_LsuL1_ABORD_lane0)) && (! execute_ctrl4_down_LsuL1_SKIP_WRITE_lane0)) && (! execute_ctrl4_down_LsuL1_MISS_lane0)) && (! execute_ctrl4_down_LsuL1_MISS_UNIQUE_lane0)) && (! execute_ctrl4_down_LsuL1_HAZARD_lane0));
  assign LsuL1TileLinkPlugin_logic_down_a_fire = (LsuL1TileLinkPlugin_logic_down_a_valid && LsuL1TileLinkPlugin_logic_down_a_ready);
  assign LsuL1TileLinkPlugin_logic_down_a_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == LsuL1TileLinkPlugin_logic_down_a_payload_opcode)) || (A_PUT_PARTIAL_DATA == LsuL1TileLinkPlugin_logic_down_a_payload_opcode))) || (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat == _zz_LsuL1TileLinkPlugin_logic_down_a_tracker_last));
  assign when_LsuL1Bus_l151 = (LsuL1TileLinkPlugin_logic_down_a_fire && LsuL1TileLinkPlugin_logic_down_a_tracker_last);
  assign LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel = (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock ? LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_selReg : LsuL1Plugin_logic_bus_read_cmd_valid);
  assign LsuL1TileLinkPlugin_logic_down_a_payload_param = 3'b000;
  assign LsuL1TileLinkPlugin_logic_down_a_payload_size = 3'b110;
  assign LsuL1TileLinkPlugin_logic_down_a_payload_mask = 8'hff;
  assign LsuL1TileLinkPlugin_logic_down_a_payload_data = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_data;
  assign LsuL1TileLinkPlugin_logic_down_a_payload_corrupt = 1'b0;
  always @(*) begin
    if(LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) begin
      LsuL1TileLinkPlugin_logic_down_a_valid = LsuL1Plugin_logic_bus_read_cmd_valid;
    end else begin
      LsuL1TileLinkPlugin_logic_down_a_valid = LsuL1Plugin_logic_bus_write_cmd_valid;
    end
  end

  always @(*) begin
    if(LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) begin
      LsuL1TileLinkPlugin_logic_down_a_payload_opcode = A_GET;
    end else begin
      LsuL1TileLinkPlugin_logic_down_a_payload_opcode = A_PUT_FULL_DATA;
    end
  end

  always @(*) begin
    if(LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) begin
      LsuL1TileLinkPlugin_logic_down_a_payload_source = 1'b0;
    end else begin
      LsuL1TileLinkPlugin_logic_down_a_payload_source = 1'b0;
    end
    LsuL1TileLinkPlugin_logic_down_a_payload_source[0] = LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel;
  end

  always @(*) begin
    if(LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) begin
      LsuL1TileLinkPlugin_logic_down_a_payload_address = LsuL1Plugin_logic_bus_read_cmd_payload_address;
    end else begin
      LsuL1TileLinkPlugin_logic_down_a_payload_address = LsuL1Plugin_logic_bus_write_cmd_payload_fragment_address;
    end
    LsuL1TileLinkPlugin_logic_down_a_payload_address[5 : 3] = LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat;
  end

  assign LsuL1Plugin_logic_bus_write_cmd_ready = ((! LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel) && LsuL1TileLinkPlugin_logic_down_a_ready);
  assign LsuL1Plugin_logic_bus_read_cmd_ready = (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel && LsuL1TileLinkPlugin_logic_down_a_ready);
  assign LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel = LsuL1TileLinkPlugin_logic_down_d_payload_source[0];
  assign LsuL1Plugin_logic_bus_read_rsp_valid = (LsuL1TileLinkPlugin_logic_down_d_valid && LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel);
  assign LsuL1Plugin_logic_bus_read_rsp_payload_data = LsuL1TileLinkPlugin_logic_down_d_payload_data;
  assign LsuL1Plugin_logic_bus_read_rsp_payload_error = (LsuL1TileLinkPlugin_logic_down_d_payload_denied || LsuL1TileLinkPlugin_logic_down_d_payload_corrupt);
  assign LsuL1Plugin_logic_bus_write_rsp_valid = (LsuL1TileLinkPlugin_logic_down_d_valid && (! LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel));
  assign LsuL1Plugin_logic_bus_write_rsp_payload_error = (LsuL1TileLinkPlugin_logic_down_d_payload_denied || LsuL1TileLinkPlugin_logic_down_d_payload_corrupt);
  assign LsuL1TileLinkPlugin_logic_down_d_ready = (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onD_sel ? LsuL1Plugin_logic_bus_read_rsp_ready : 1'b1);
  assign PcPlugin_logic_forcedSpawn = (|{TrapPlugin_logic_harts_0_trap_pcPort_valid,{early0_BranchPlugin_logic_pcPort_valid,BtbPlugin_logic_pcPort_valid}});
  assign PcPlugin_logic_harts_0_self_pc = (PcPlugin_logic_harts_0_self_state + _zz_PcPlugin_logic_harts_0_self_pc);
  assign PcPlugin_logic_harts_0_self_flow_valid = 1'b1;
  assign PcPlugin_logic_harts_0_self_flow_payload_fault = PcPlugin_logic_harts_0_self_fault;
  assign PcPlugin_logic_harts_0_self_flow_payload_pc = PcPlugin_logic_harts_0_self_pc;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid = 1'b1;
  assign PcPlugin_logic_harts_0_aggregator_valids_0 = ((TrapPlugin_logic_harts_0_trap_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_0_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_1 = ((early0_BranchPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_1_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_2 = ((BtbPlugin_logic_pcPort_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_2_laneValid);
  assign PcPlugin_logic_harts_0_aggregator_valids_3 = ((PcPlugin_logic_harts_0_self_flow_valid && 1'b1) && PcPlugin_logic_harts_0_aggregator_sortedByPriority_3_laneValid);
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh = {PcPlugin_logic_harts_0_aggregator_valids_3,{PcPlugin_logic_harts_0_aggregator_valids_2,{PcPlugin_logic_harts_0_aggregator_valids_1,PcPlugin_logic_harts_0_aggregator_valids_0}}};
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_1 = _zz_PcPlugin_logic_harts_0_aggregator_oh[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_2 = _zz_PcPlugin_logic_harts_0_aggregator_oh[1];
  assign _zz_PcPlugin_logic_harts_0_aggregator_oh_3 = _zz_PcPlugin_logic_harts_0_aggregator_oh[2];
  always @(*) begin
    _zz_PcPlugin_logic_harts_0_aggregator_oh_4[0] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_1 && (! 1'b0));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_4[1] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_2 && (! _zz_PcPlugin_logic_harts_0_aggregator_oh_1));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_4[2] = (_zz_PcPlugin_logic_harts_0_aggregator_oh_3 && (! (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1})));
    _zz_PcPlugin_logic_harts_0_aggregator_oh_4[3] = (_zz_PcPlugin_logic_harts_0_aggregator_oh[3] && (! (|{_zz_PcPlugin_logic_harts_0_aggregator_oh_3,{_zz_PcPlugin_logic_harts_0_aggregator_oh_2,_zz_PcPlugin_logic_harts_0_aggregator_oh_1}})));
  end

  assign PcPlugin_logic_harts_0_aggregator_oh = _zz_PcPlugin_logic_harts_0_aggregator_oh_4;
  assign _zz_PcPlugin_logic_harts_0_aggregator_target = PcPlugin_logic_harts_0_aggregator_oh[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_1 = PcPlugin_logic_harts_0_aggregator_oh[1];
  assign _zz_PcPlugin_logic_harts_0_aggregator_target_2 = PcPlugin_logic_harts_0_aggregator_oh[3];
  assign PcPlugin_logic_harts_0_aggregator_target = (((_zz_PcPlugin_logic_harts_0_aggregator_target ? TrapPlugin_logic_harts_0_trap_pcPort_payload_pc : 32'h0) | (_zz_PcPlugin_logic_harts_0_aggregator_target_1 ? early0_BranchPlugin_logic_pcPort_payload_pc : 32'h0)) | (_zz_PcPlugin_logic_harts_0_aggregator_target_2 ? PcPlugin_logic_harts_0_self_flow_payload_pc : 32'h0));
  assign PcPlugin_logic_harts_0_aggregator_fault = _zz_PcPlugin_logic_harts_0_aggregator_fault[0];
  assign _zz_PcPlugin_logic_harts_0_aggregator_fault_1 = PcPlugin_logic_harts_0_aggregator_oh[2];
  assign when_PcPlugin_l80 = (|_zz_PcPlugin_logic_harts_0_aggregator_fault_1);
  assign PcPlugin_logic_harts_0_holdComb = (|TrapPlugin_logic_harts_0_trap_fsm_holdPort);
  assign PcPlugin_logic_harts_0_output_valid = (! PcPlugin_logic_harts_0_holdReg);
  assign PcPlugin_logic_harts_0_output_payload_fault = PcPlugin_logic_harts_0_aggregator_fault_1;
  always @(*) begin
    PcPlugin_logic_harts_0_output_payload_pc = PcPlugin_logic_harts_0_aggregator_target_1;
    PcPlugin_logic_harts_0_output_payload_pc[1 : 0] = 2'b00;
  end

  assign PcPlugin_logic_harts_0_output_fire = (PcPlugin_logic_harts_0_output_valid && PcPlugin_logic_harts_0_output_ready);
  assign fetch_logic_ctrls_0_up_valid = PcPlugin_logic_harts_0_output_valid;
  assign PcPlugin_logic_harts_0_output_ready = fetch_logic_ctrls_0_up_ready;
  assign fetch_logic_ctrls_0_up_Fetch_WORD_PC = PcPlugin_logic_harts_0_output_payload_pc;
  assign fetch_logic_ctrls_0_up_Fetch_PC_FAULT = PcPlugin_logic_harts_0_output_payload_fault;
  always @(*) begin
    fetch_logic_ctrls_0_up_Fetch_ID = 10'bxxxxxxxxxx;
    fetch_logic_ctrls_0_up_Fetch_ID = PcPlugin_logic_harts_0_self_id;
  end

  assign PcPlugin_logic_holdHalter_doIt = PcPlugin_logic_harts_0_holdComb;
  assign fetch_logic_ctrls_0_haltRequest_PcPlugin_l133 = PcPlugin_logic_holdHalter_doIt;
  always @(*) begin
    HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_value;
    if(HistoryPlugin_logic_onFetch_ports_0_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_0_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_1_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_1_payload_history;
    end
    if(HistoryPlugin_logic_onFetch_ports_2_valid) begin
      HistoryPlugin_logic_onFetch_valueNext = HistoryPlugin_logic_onFetch_ports_2_payload_history;
    end
  end

  assign HistoryPlugin_logic_onFetch_ports_0_valid = (|BtbPlugin_logic_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_0_payload_history = BtbPlugin_logic_historyPort_payload_history;
  assign HistoryPlugin_logic_onFetch_ports_1_valid = (|early0_BranchPlugin_logic_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_1_payload_history = early0_BranchPlugin_logic_historyPort_payload_history;
  assign HistoryPlugin_logic_onFetch_ports_2_valid = (|TrapPlugin_logic_harts_0_trap_historyPort_valid);
  assign HistoryPlugin_logic_onFetch_ports_2_payload_history = TrapPlugin_logic_harts_0_trap_historyPort_payload_history;
  assign fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY = HistoryPlugin_logic_onFetch_valueNext;
  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = 2'b00;
    if(!when_MmuPlugin_l512) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = 2'b11;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = (MmuPlugin_logic_refill_storageOhReg[0] ? _zz_FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask : 2'b00);
            if(when_MmuPlugin_l455) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask = 2'b00;
            end
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address = 5'bxxxxx;
    if(!when_MmuPlugin_l512) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[16 : 12];
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l512) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = 15'bxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 17];
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value == 1'b1);
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflow = (FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc && FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext = (FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value + FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
    if(FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_willClear) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext = 1'b0;
    end
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
    if(!when_MmuPlugin_l512) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b1;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = (MmuPlugin_logic_refill_storageOhReg[0] ? 1'b1 : 1'b0);
              if(when_MmuPlugin_l455_2) begin
                FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = 5'bxxxxx;
    if(!when_MmuPlugin_l512) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[26 : 22];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l512) begin
      FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = 5'bxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 27];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = 10'bxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd22);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc = 1'b1;
  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflow = (FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc && FetchL1Plugin_logic_translationStorage_logic_sl_1_allocId_willIncrement);
  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = 3'b000;
    if(!when_MmuPlugin_l512) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = 3'b111;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = _zz_LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[2:0];
            if(when_MmuPlugin_l455_1) begin
              LsuPlugin_logic_translationStorage_logic_sl_0_write_mask = 3'b000;
            end
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_address = 5'bxxxxx;
    if(!when_MmuPlugin_l512) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_address = MmuPlugin_logic_refill_virtual[16 : 12];
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l512) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = 15'bxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 17];
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = 20'bxxxxxxxxxxxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 >>> 4'd12);
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement = 1'b1;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willClear = 1'b0;
  assign LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc = (LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value == 2'b10);
  assign LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflow = (LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflowIfInc && LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willIncrement);
  always @(*) begin
    if(LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willOverflow) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = 2'b00;
    end else begin
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = (LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value + _zz_LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext);
    end
    if(LsuPlugin_logic_translationStorage_logic_sl_0_allocId_willClear) begin
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext = 2'b00;
    end
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
    if(!when_MmuPlugin_l512) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b1;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = (MmuPlugin_logic_refill_storageOhReg[1] ? 1'b1 : 1'b0);
              if(when_MmuPlugin_l455_3) begin
                LsuPlugin_logic_translationStorage_logic_sl_1_write_mask = 1'b0;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_address = 5'bxxxxx;
    if(!when_MmuPlugin_l512) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_invalidate_counter;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_address = MmuPlugin_logic_refill_virtual[26 : 22];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'bx;
    if(!when_MmuPlugin_l512) begin
      LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b0;
    end
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = 5'bxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress = MmuPlugin_logic_refill_virtual[31 : 27];
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = 10'bxxxxxxxxxx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress = (MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 >>> 5'd22);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead = MmuPlugin_logic_refill_load_flags_R;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite = (MmuPlugin_logic_refill_load_flags_W && MmuPlugin_logic_refill_load_flags_D);
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute = MmuPlugin_logic_refill_load_flags_X;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser = MmuPlugin_logic_refill_load_flags_U;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement = 1'b1;
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willClear = 1'b0;
  assign LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc = 1'b1;
  assign LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflow = (LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willOverflowIfInc && LsuPlugin_logic_translationStorage_logic_sl_1_allocId_willIncrement);
  assign MmuPlugin_logic_isMachine = (PrivilegedPlugin_logic_harts_0_privilege == 2'b11);
  assign MmuPlugin_logic_isSupervisor = (PrivilegedPlugin_logic_harts_0_privilege == 2'b01);
  assign MmuPlugin_logic_isUser = (PrivilegedPlugin_logic_harts_0_privilege == 2'b00);
  always @(*) begin
    MmuPlugin_api_fetchTranslationEnable = (MmuPlugin_logic_satp_mode == 1'b1);
    if(MmuPlugin_logic_isMachine) begin
      MmuPlugin_api_fetchTranslationEnable = 1'b0;
    end
  end

  always @(*) begin
    MmuPlugin_api_lsuTranslationEnable = (MmuPlugin_logic_satp_mode == 1'b1);
    if(when_MmuPlugin_l275) begin
      MmuPlugin_api_lsuTranslationEnable = 1'b0;
    end
    if(MmuPlugin_logic_isMachine) begin
      if(when_MmuPlugin_l277) begin
        MmuPlugin_api_lsuTranslationEnable = 1'b0;
      end
    end
  end

  assign when_MmuPlugin_l275 = ((! PrivilegedPlugin_logic_harts_0_m_status_mprv) && MmuPlugin_logic_isMachine);
  assign when_MmuPlugin_l277 = ((! PrivilegedPlugin_logic_harts_0_m_status_mprv) || (PrivilegedPlugin_logic_harts_0_m_status_mpp == 2'b11));
  assign LsuPlugin_logic_onAddress0_translationPort_logic_read_0_readAddress = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[16 : 12];
  assign _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid = LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_rd_data;
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[0];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_virtualAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[15 : 1];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_physicalAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[35 : 16];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowRead = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[36];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowWrite = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[37];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowExecute = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[38];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowUser = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid[39];
  always @(*) begin
    execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0[0] = (execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_virtualAddress == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[31 : 17]);
    execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0[1] = (execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_virtualAddress == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[31 : 17]);
    execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0[2] = (execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_virtualAddress == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[31 : 17]);
  end

  always @(*) begin
    execute_ctrl3_down_MMU_L0_HITS_lane0[0] = (execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[0] && execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid);
    execute_ctrl3_down_MMU_L0_HITS_lane0[1] = (execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[1] && execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid);
    execute_ctrl3_down_MMU_L0_HITS_lane0[2] = (execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0[2] && execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_valid);
  end

  assign _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid = LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_rd_data;
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[0];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_virtualAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[15 : 1];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_physicalAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[35 : 16];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowRead = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[36];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowWrite = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[37];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowExecute = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[38];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowUser = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid[39];
  assign _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid = LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_rd_data;
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[0];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_virtualAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[15 : 1];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_physicalAddress = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[35 : 16];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowRead = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[36];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowWrite = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[37];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowExecute = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[38];
  assign execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowUser = _zz_execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid[39];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_read_1_readAddress = execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[26 : 22];
  assign _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid = LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_rd_data;
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[0];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_virtualAddress = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[5 : 1];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_physicalAddress = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[15 : 6];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowRead = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[16];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowWrite = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[17];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowExecute = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[18];
  assign execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowUser = _zz_execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid[19];
  assign execute_ctrl2_down_MMU_L1_HITS_PRE_VALID_lane0[0] = (execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_virtualAddress == execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0[31 : 27]);
  assign execute_ctrl3_down_MMU_L1_HITS_lane0[0] = (execute_ctrl3_down_MMU_L1_HITS_PRE_VALID_lane0[0] && execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid);
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits = {execute_ctrl3_down_MMU_L1_HITS_lane0,execute_ctrl3_down_MMU_L0_HITS_lane0};
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hit = (|LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits);
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits;
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[1];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[2];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_3 = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0[3];
  always @(*) begin
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[0] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[1] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1 && (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0));
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[2] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2 && (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_1));
    _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[3] = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_3 && (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_2));
  end

  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_1 = (|{LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1,LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0});
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_range_0_to_2 = (|{LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_2,{LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_1,LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hits_bools_0}});
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[0];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[1];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[2];
  assign _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh[3];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_4[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser = _zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser[0];
  assign LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated = (((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute ? {_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_1} : 32'h0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_1 ? {_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_2,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_3} : 32'h0)) | ((_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_2 ? {_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_4,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_5} : 32'h0) | (_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute_3 ? {_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_6,_zz_LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated_7} : 32'h0)));
  always @(*) begin
    LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup = MmuPlugin_api_lsuTranslationEnable;
    if(execute_ctrl3_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0) begin
      LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_HAZARD_lane0 = 1'b0;
    end else begin
      execute_ctrl3_down_MMU_HAZARD_lane0 = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_REFILL_lane0 = (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_hit);
    end else begin
      execute_ctrl3_down_MMU_REFILL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_TRANSLATED_lane0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineTranslated;
    end else begin
      execute_ctrl3_down_MMU_TRANSLATED_lane0 = execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0 = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute && (! (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor)));
    end else begin
      execute_ctrl3_down_MMU_ALLOW_EXECUTE_lane0 = 1'b1;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_ALLOW_READ_lane0 = (LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      execute_ctrl3_down_MMU_ALLOW_READ_lane0 = 1'b1;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_ALLOW_WRITE_lane0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      execute_ctrl3_down_MMU_ALLOW_WRITE_lane0 = 1'b1;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_PAGE_FAULT_lane0 = (((LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor) && (! MmuPlugin_logic_status_sum)) || ((! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_lineAllowUser) && MmuPlugin_logic_isUser));
    end else begin
      execute_ctrl3_down_MMU_PAGE_FAULT_lane0 = 1'b0;
    end
  end

  always @(*) begin
    if(LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup) begin
      execute_ctrl3_down_MMU_ACCESS_FAULT_lane0 = 1'b0;
    end else begin
      execute_ctrl3_down_MMU_ACCESS_FAULT_lane0 = 1'b0;
    end
  end

  assign execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0 = (! LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_requireMmuLockup);
  assign execute_ctrl3_down_MMU_WAYS_OH_lane0 = LsuPlugin_logic_onAddress0_translationPort_logic_ctrl_oh;
  assign execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_0 = {execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress,execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0]};
  assign execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_1 = {execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress,execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0]};
  assign execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_2 = {execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_physicalAddress,execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[11 : 0]};
  assign execute_ctrl3_down_MMU_WAYS_PHYSICAL_lane0_3 = {execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress,execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0[21 : 0]};
  assign FetchL1Plugin_logic_translationPort_logic_read_0_readAddress = fetch_logic_ctrls_1_down_Fetch_WORD_PC[16 : 12];
  assign _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_rd_data;
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[0];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_virtualAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[15 : 1];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[35 : 16];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowRead = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[36];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowWrite = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[37];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowExecute = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[38];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_allowUser = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid[39];
  always @(*) begin
    fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[0] = (fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_virtualAddress == fetch_logic_ctrls_1_down_Fetch_WORD_PC[31 : 17]);
    fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[1] = (fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_virtualAddress == fetch_logic_ctrls_1_down_Fetch_WORD_PC[31 : 17]);
  end

  always @(*) begin
    fetch_logic_ctrls_1_down_MMU_L0_HITS[0] = (fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[0] && fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_valid);
    fetch_logic_ctrls_1_down_MMU_L0_HITS[1] = (fetch_logic_ctrls_1_down_MMU_L0_HITS_PRE_VALID[1] && fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid);
  end

  assign _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid = FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_rd_data;
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[0];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_virtualAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[15 : 1];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[35 : 16];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowRead = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[36];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowWrite = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[37];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowExecute = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[38];
  assign fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_allowUser = _zz_fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_valid[39];
  assign FetchL1Plugin_logic_translationPort_logic_read_1_readAddress = fetch_logic_ctrls_1_down_Fetch_WORD_PC[26 : 22];
  assign _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid = FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_rd_data;
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[0];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_virtualAddress = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[5 : 1];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[15 : 6];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowRead = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[16];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowWrite = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[17];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowExecute = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[18];
  assign fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_allowUser = _zz_fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid[19];
  assign fetch_logic_ctrls_1_down_MMU_L1_HITS_PRE_VALID[0] = (fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_virtualAddress == fetch_logic_ctrls_1_down_Fetch_WORD_PC[31 : 27]);
  assign fetch_logic_ctrls_1_down_MMU_L1_HITS[0] = (fetch_logic_ctrls_1_down_MMU_L1_HITS_PRE_VALID[0] && fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_valid);
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits = {fetch_logic_ctrls_1_down_MMU_L1_HITS,fetch_logic_ctrls_1_down_MMU_L0_HITS};
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hit = (|FetchL1Plugin_logic_translationPort_logic_ctrl_hits);
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0 = FetchL1Plugin_logic_translationPort_logic_ctrl_hits;
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0 = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1 = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0[1];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_2 = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0[2];
  always @(*) begin
    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh[0] = (FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0 && (! 1'b0));
    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh[1] = (FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1 && (! FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0));
    _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh[2] = (FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_2 && (! FetchL1Plugin_logic_translationPort_logic_ctrl_hits_range_0_to_1));
  end

  assign FetchL1Plugin_logic_translationPort_logic_ctrl_hits_range_0_to_1 = (|{FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_1,FetchL1Plugin_logic_translationPort_logic_ctrl_hits_bools_0});
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_oh = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute = FetchL1Plugin_logic_translationPort_logic_ctrl_oh[0];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 = FetchL1Plugin_logic_translationPort_logic_ctrl_oh[1];
  assign _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 = FetchL1Plugin_logic_translationPort_logic_ctrl_oh[2];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_3[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser = _zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser[0];
  assign FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated = (((_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute ? {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress,_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated} : 32'h0) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_1 ? {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress,_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated_1} : 32'h0)) | (_zz_FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute_2 ? {fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[21 : 0]} : 32'h0));
  always @(*) begin
    FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup = MmuPlugin_api_fetchTranslationEnable;
    if(_zz_1) begin
      FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_HAZARD = 1'b0;
    end else begin
      fetch_logic_ctrls_1_down_MMU_HAZARD = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_REFILL = (! FetchL1Plugin_logic_translationPort_logic_ctrl_hit);
    end else begin
      fetch_logic_ctrls_1_down_MMU_REFILL = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_TRANSLATED = FetchL1Plugin_logic_translationPort_logic_ctrl_lineTranslated;
    end else begin
      fetch_logic_ctrls_1_down_MMU_TRANSLATED = fetch_logic_ctrls_1_down_Fetch_WORD_PC;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE = (FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute && (! (FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor)));
    end else begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE = 1'b1;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_READ = (FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowRead || (MmuPlugin_logic_status_mxr && FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowExecute));
    end else begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_READ = 1'b1;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE = FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowWrite;
    end else begin
      fetch_logic_ctrls_1_down_MMU_ALLOW_WRITE = 1'b1;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_PAGE_FAULT = (((FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser && MmuPlugin_logic_isSupervisor) && (! MmuPlugin_logic_status_sum)) || ((! FetchL1Plugin_logic_translationPort_logic_ctrl_lineAllowUser) && MmuPlugin_logic_isUser));
    end else begin
      fetch_logic_ctrls_1_down_MMU_PAGE_FAULT = 1'b0;
    end
  end

  always @(*) begin
    if(FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup) begin
      fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT = 1'b0;
    end else begin
      fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT = 1'b0;
    end
  end

  assign fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION = (! FetchL1Plugin_logic_translationPort_logic_ctrl_requireMmuLockup);
  assign fetch_logic_ctrls_1_down_MMU_WAYS_OH = FetchL1Plugin_logic_translationPort_logic_ctrl_oh;
  assign fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_0 = {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_0_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0]};
  assign fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_1 = {fetch_logic_ctrls_1_down_MMU_L0_ENTRIES_1_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[11 : 0]};
  assign fetch_logic_ctrls_1_down_MMU_WAYS_PHYSICAL_2 = {fetch_logic_ctrls_1_down_MMU_L1_ENTRIES_0_physicalAddress,fetch_logic_ctrls_1_down_Fetch_WORD_PC[21 : 0]};
  assign MmuPlugin_logic_refill_wantExit = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_wantStart = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
        MmuPlugin_logic_refill_wantStart = 1'b1;
      end
    endcase
  end

  assign MmuPlugin_logic_refill_wantKill = 1'b0;
  assign MmuPlugin_logic_refill_busy = (! (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_IDLE));
  always @(*) begin
    MmuPlugin_logic_refill_cacheRefillAnySet = 1'b0;
    if(when_MmuPlugin_l395) begin
      MmuPlugin_logic_refill_cacheRefillAnySet = MmuPlugin_logic_accessBus_rsp_payload_waitAny;
    end
  end

  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_ready = MmuPlugin_logic_refill_arbiter_io_inputs_0_ready;
  always @(*) begin
    MmuPlugin_logic_refill_arbiter_io_output_ready = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
        if(MmuPlugin_logic_refill_arbiter_io_output_valid) begin
          MmuPlugin_logic_refill_arbiter_io_output_ready = 1'b1;
        end
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_events_onStorage_0_waiting = (MmuPlugin_logic_refill_busy && MmuPlugin_logic_refill_storageOhReg[0]);
  assign MmuPlugin_logic_refill_events_onStorage_1_waiting = (MmuPlugin_logic_refill_busy && MmuPlugin_logic_refill_storageOhReg[1]);
  assign MmuPlugin_logic_refill_load_readed = MmuPlugin_logic_refill_load_rsp_payload_data[31 : 0];
  assign when_MmuPlugin_l395 = (MmuPlugin_logic_accessBus_rsp_valid && MmuPlugin_logic_accessBus_rsp_payload_redo);
  always @(*) begin
    MmuPlugin_logic_accessBus_cmd_valid = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
        if(when_MmuPlugin_l470) begin
          MmuPlugin_logic_accessBus_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_CMD_1 : begin
        if(when_MmuPlugin_l470_1) begin
          MmuPlugin_logic_accessBus_cmd_valid = 1'b1;
        end
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_accessBus_cmd_payload_address = MmuPlugin_logic_refill_load_address;
  assign MmuPlugin_logic_accessBus_cmd_payload_size = 2'b10;
  assign _zz_MmuPlugin_logic_refill_load_flags_V = MmuPlugin_logic_refill_load_readed;
  assign MmuPlugin_logic_refill_load_flags_V = _zz_MmuPlugin_logic_refill_load_flags_V[0];
  assign MmuPlugin_logic_refill_load_flags_R = _zz_MmuPlugin_logic_refill_load_flags_V[1];
  assign MmuPlugin_logic_refill_load_flags_W = _zz_MmuPlugin_logic_refill_load_flags_V[2];
  assign MmuPlugin_logic_refill_load_flags_X = _zz_MmuPlugin_logic_refill_load_flags_V[3];
  assign MmuPlugin_logic_refill_load_flags_U = _zz_MmuPlugin_logic_refill_load_flags_V[4];
  assign MmuPlugin_logic_refill_load_flags_G = _zz_MmuPlugin_logic_refill_load_flags_V[5];
  assign MmuPlugin_logic_refill_load_flags_A = _zz_MmuPlugin_logic_refill_load_flags_V[6];
  assign MmuPlugin_logic_refill_load_flags_D = _zz_MmuPlugin_logic_refill_load_flags_V[7];
  assign MmuPlugin_logic_refill_load_leaf = (MmuPlugin_logic_refill_load_flags_R || MmuPlugin_logic_refill_load_flags_X);
  assign MmuPlugin_logic_refill_load_reservedFault = (|(MmuPlugin_logic_refill_load_readed & 32'h0));
  always @(*) begin
    MmuPlugin_logic_refill_load_exception = (((((! MmuPlugin_logic_refill_load_flags_V) || ((! MmuPlugin_logic_refill_load_flags_R) && MmuPlugin_logic_refill_load_flags_W)) || MmuPlugin_logic_refill_load_rsp_payload_error) || ((! MmuPlugin_logic_refill_load_leaf) && ((MmuPlugin_logic_refill_load_flags_D || MmuPlugin_logic_refill_load_flags_A) || MmuPlugin_logic_refill_load_flags_U))) || MmuPlugin_logic_refill_load_reservedFault);
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(when_MmuPlugin_l479) begin
          MmuPlugin_logic_refill_load_exception = 1'b1;
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_load_levelException_0 = 1'b0;
  always @(*) begin
    MmuPlugin_logic_refill_load_levelException_1 = 1'b0;
    if(when_MmuPlugin_l416) begin
      MmuPlugin_logic_refill_load_levelException_1 = 1'b1;
    end
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_nextLevelBase = 32'h0;
    MmuPlugin_logic_refill_load_nextLevelBase[21 : 12] = MmuPlugin_logic_refill_load_readed[19 : 10];
    MmuPlugin_logic_refill_load_nextLevelBase[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0 = 32'h0;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[21 : 12] = MmuPlugin_logic_refill_load_readed[19 : 10];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_0[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  always @(*) begin
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1 = 32'h0;
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[21 : 12] = MmuPlugin_logic_refill_virtual[21 : 12];
    MmuPlugin_logic_refill_load_levelToPhysicalAddress_1[31 : 22] = MmuPlugin_logic_refill_load_readed[29 : 20];
  end

  assign when_MmuPlugin_l416 = (MmuPlugin_logic_refill_load_readed[19 : 10] != 10'h0);
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b0;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(_zz_57) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
            end
            if(_zz_57) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
            end
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              if(_zz_57) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
              end
              if(_zz_57) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid = 1'b1;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(_zz_57) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = MmuPlugin_logic_refill_fetch_0_pageFault;
            end
            if(_zz_57) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = MmuPlugin_logic_refill_fetch_0_pageFault;
            end
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              if(_zz_57) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = MmuPlugin_logic_refill_fetch_1_pageFault;
              end
              if(_zz_57) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault = MmuPlugin_logic_refill_fetch_1_pageFault;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = 1'bx;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(_zz_57) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = MmuPlugin_logic_refill_fetch_0_accessFault;
            end
            if(_zz_57) begin
              TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = MmuPlugin_logic_refill_fetch_0_accessFault;
            end
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(when_MmuPlugin_l487) begin
              if(_zz_57) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = MmuPlugin_logic_refill_fetch_1_accessFault;
              end
              if(_zz_57) begin
                TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault = MmuPlugin_logic_refill_fetch_1_accessFault;
              end
            end
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign MmuPlugin_logic_refill_fetch_0_pteFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_0) || (! MmuPlugin_logic_refill_load_flags_A));
  assign MmuPlugin_logic_refill_fetch_0_leafAccessFault = 1'b0;
  assign MmuPlugin_logic_refill_fetch_0_pageFault = ((! MmuPlugin_logic_refill_load_rsp_payload_error) && MmuPlugin_logic_refill_fetch_0_pteFault);
  assign MmuPlugin_logic_refill_fetch_0_accessFault = (MmuPlugin_logic_refill_load_rsp_payload_error || ((! MmuPlugin_logic_refill_fetch_0_pteFault) && MmuPlugin_logic_refill_fetch_0_leafAccessFault));
  assign MmuPlugin_logic_refill_fetch_1_pteFault = ((MmuPlugin_logic_refill_load_exception || MmuPlugin_logic_refill_load_levelException_1) || (! MmuPlugin_logic_refill_load_flags_A));
  assign MmuPlugin_logic_refill_fetch_1_leafAccessFault = 1'b0;
  assign MmuPlugin_logic_refill_fetch_1_pageFault = ((! MmuPlugin_logic_refill_load_rsp_payload_error) && MmuPlugin_logic_refill_fetch_1_pteFault);
  assign MmuPlugin_logic_refill_fetch_1_accessFault = (MmuPlugin_logic_refill_load_rsp_payload_error || ((! MmuPlugin_logic_refill_fetch_1_pteFault) && MmuPlugin_logic_refill_fetch_1_leafAccessFault));
  assign TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready = MmuPlugin_logic_invalidate_arbiter_io_inputs_0_ready;
  always @(*) begin
    MmuPlugin_logic_invalidate_arbiter_io_output_ready = 1'b0;
    if(!when_MmuPlugin_l512) begin
      if(when_MmuPlugin_l526) begin
        MmuPlugin_logic_invalidate_arbiter_io_output_ready = 1'b1;
      end
    end
  end

  assign when_MmuPlugin_l512 = (! MmuPlugin_logic_invalidate_busy);
  assign when_MmuPlugin_l526 = (&MmuPlugin_logic_invalidate_counter);
  assign PmpPlugin_logic_isMachine = (PrivilegedPlugin_logic_harts_0_privilege == 2'b11);
  assign PmpPlugin_logic_instructionShouldHit = (! PmpPlugin_logic_isMachine);
  assign PmpPlugin_logic_dataShouldHit = ((! PmpPlugin_logic_isMachine) || (PrivilegedPlugin_logic_harts_0_m_status_mprv && (PrivilegedPlugin_logic_harts_0_m_status_mpp != 2'b11)));
  assign FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort = (PmpPlugin_logic_dataShouldHit || 1'b0);
  assign FetchL1Plugin_logic_pmpPort_logic_torCmpAddress = (fetch_logic_ctrls_1_down_MMU_TRANSLATED >>> 4'd12);
  assign fetch_logic_ctrls_0_down_FetchL1Plugin_logic_pmpPort_logic_NEED_HIT = ((PmpPlugin_logic_instructionShouldHit && 1'b1) || (FetchL1Plugin_logic_pmpPort_logic_dataShouldHitPort && (1'b0 || 1'b0)));
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_pmpPort_ACCESS_FAULT = 1'b0;
  assign LsuPlugin_logic_pmpPort_logic_dataShouldHitPort = (PmpPlugin_logic_dataShouldHit || execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0);
  assign LsuPlugin_logic_pmpPort_logic_torCmpAddress = (execute_ctrl3_down_MMU_TRANSLATED_lane0 >>> 4'd12);
  assign execute_ctrl2_down_LsuPlugin_logic_pmpPort_logic_NEED_HIT_lane0 = ((PmpPlugin_logic_instructionShouldHit && 1'b0) || (LsuPlugin_logic_pmpPort_logic_dataShouldHitPort && (execute_ctrl2_down_LsuL1_LOAD_lane0 || execute_ctrl2_down_LsuL1_STORE_lane0)));
  assign execute_ctrl4_down_LsuPlugin_logic_pmpPort_ACCESS_FAULT_lane0 = 1'b0;
  assign LsuTileLinkPlugin_logic_bridge_cmdHash = LsuPlugin_logic_bus_cmd_payload_address[9 : 2];
  assign LsuTileLinkPlugin_logic_bridge_down_a_valid = LsuPlugin_logic_bus_cmd_valid;
  assign LsuPlugin_logic_bus_cmd_ready = LsuTileLinkPlugin_logic_bridge_down_a_ready;
  assign _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode = (LsuPlugin_logic_bus_cmd_payload_write ? A_PUT_FULL_DATA : A_GET);
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode = _zz_LsuTileLinkPlugin_logic_bridge_down_a_payload_opcode;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_param = 3'b000;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_address = LsuPlugin_logic_bus_cmd_payload_address;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_size = LsuPlugin_logic_bus_cmd_payload_size;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_mask = LsuPlugin_logic_bus_cmd_payload_mask;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_data = LsuPlugin_logic_bus_cmd_payload_data;
  assign LsuTileLinkPlugin_logic_bridge_down_a_payload_corrupt = 1'b0;
  assign LsuTileLinkPlugin_logic_bridge_down_d_ready = 1'b1;
  assign LsuPlugin_logic_bus_rsp_valid = LsuTileLinkPlugin_logic_bridge_down_d_valid;
  assign LsuPlugin_logic_bus_rsp_payload_error = LsuTileLinkPlugin_logic_bridge_down_d_payload_denied;
  assign LsuPlugin_logic_bus_rsp_payload_data = LsuTileLinkPlugin_logic_bridge_down_d_payload_data;
  assign fetch_logic_flushes_0_doIt = (|{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),{(LsuPlugin_logic_flushPort_valid && 1'b1),((BtbPlugin_logic_flushPort_valid && _zz_fetch_logic_flushes_0_doIt) && (_zz_fetch_logic_flushes_0_doIt_1 || _zz_fetch_logic_flushes_0_doIt_2))}}}}});
  assign fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48 = fetch_logic_flushes_0_doIt;
  assign fetch_logic_flushes_1_doIt = (|{(DecoderPlugin_logic_laneLogic_0_flushPort_valid && 1'b1),{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}}});
  assign fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l50 = fetch_logic_flushes_1_doIt;
  assign PerformanceCounterPlugin_logic_events_sums_0 = _zz_PerformanceCounterPlugin_logic_events_sums_0_1;
  assign PerformanceCounterPlugin_logic_events_sums_1 = _zz_PerformanceCounterPlugin_logic_events_sums_1_1;
  assign PerformanceCounterPlugin_logic_events_sums_2 = _zz_PerformanceCounterPlugin_logic_events_sums_2_1;
  assign PerformanceCounterPlugin_logic_events_sums_3 = _zz_PerformanceCounterPlugin_logic_events_sums_3_1;
  assign PerformanceCounterPlugin_logic_events_sums_4 = _zz_PerformanceCounterPlugin_logic_events_sums_4_1;
  assign PerformanceCounterPlugin_logic_events_sums_5 = _zz_PerformanceCounterPlugin_logic_events_sums_5_1;
  assign PerformanceCounterPlugin_logic_events_sums_6 = _zz_PerformanceCounterPlugin_logic_events_sums_6_1;
  assign PerformanceCounterPlugin_logic_events_sums_7 = _zz_PerformanceCounterPlugin_logic_events_sums_7_1;
  assign PerformanceCounterPlugin_logic_events_sums_8 = _zz_PerformanceCounterPlugin_logic_events_sums_8_1;
  assign PerformanceCounterPlugin_logic_events_sums_9 = _zz_PerformanceCounterPlugin_logic_events_sums_9_1;
  assign PerformanceCounterPlugin_logic_events_sums_10 = _zz_PerformanceCounterPlugin_logic_events_sums_10_1;
  assign PerformanceCounterPlugin_logic_events_sums_11 = _zz_PerformanceCounterPlugin_logic_events_sums_11_1;
  assign PerformanceCounterPlugin_logic_events_sums_12 = _zz_PerformanceCounterPlugin_logic_events_sums_12_1;
  assign PerformanceCounterPlugin_logic_events_sums_13 = _zz_PerformanceCounterPlugin_logic_events_sums_13_1;
  assign PerformanceCounterPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_wantStart = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
        PerformanceCounterPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_fsm_wantKill = 1'b0;
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        if(!PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid) begin
          if(!PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
            if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
              PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready = 1'b1;
            end
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_flusherCmd_ready = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        if(!PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid) begin
          if(PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
            PerformanceCounterPlugin_logic_fsm_flusherCmd_ready = 1'b1;
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
        PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign _zz_PerformanceCounterPlugin_logic_fsm_cmd_address = PerformanceCounterPlugin_logic_fsm_cmd_oh[0];
  assign _zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1 = PerformanceCounterPlugin_logic_fsm_cmd_oh[1];
  assign PerformanceCounterPlugin_logic_fsm_cmd_address = ((_zz_PerformanceCounterPlugin_logic_fsm_cmd_address ? 3'b001 : 3'b000) | (_zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1 ? 3'b000 : 3'b000));
  always @(*) begin
    PerformanceCounterPlugin_logic_readPort_valid = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
        PerformanceCounterPlugin_logic_readPort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
        PerformanceCounterPlugin_logic_readPort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_readPort_address = {PerformanceCounterPlugin_logic_fsm_cmd_address,PerformanceCounterPlugin_logic_fsm_carry};
  always @(*) begin
    PerformanceCounterPlugin_logic_writePort_valid = 1'b0;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
        PerformanceCounterPlugin_logic_writePort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
        PerformanceCounterPlugin_logic_writePort_valid = 1'b1;
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_writePort_address = PerformanceCounterPlugin_logic_readPort_address;
  always @(*) begin
    PerformanceCounterPlugin_logic_writePort_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
        PerformanceCounterPlugin_logic_writePort_data = _zz_PerformanceCounterPlugin_logic_writePort_data[31:0];
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
        PerformanceCounterPlugin_logic_writePort_data = _zz_PerformanceCounterPlugin_logic_writePort_data_1[31:0];
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_fsm_calc_a = (PerformanceCounterPlugin_logic_fsm_carry ? PerformanceCounterPlugin_logic_fsm_ramReaded : {PerformanceCounterPlugin_logic_fsm_ramReaded[31 : 7],_zz_PerformanceCounterPlugin_logic_fsm_calc_a});
  assign PerformanceCounterPlugin_logic_fsm_calc_b = (PerformanceCounterPlugin_logic_fsm_carry ? 8'h01 : _zz_PerformanceCounterPlugin_logic_fsm_calc_b);
  assign PerformanceCounterPlugin_logic_fsm_calc_sum = ({1'b0,PerformanceCounterPlugin_logic_fsm_calc_a} + _zz_PerformanceCounterPlugin_logic_fsm_calc_sum);
  assign PerformanceCounterPlugin_logic_fsm_idleCsrAddress = (PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid ? PerformanceCounterPlugin_logic_fsm_csrReadCmd_payload_address : PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address);
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_holdCsrWrite = 1'b1;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        PerformanceCounterPlugin_logic_fsm_holdCsrWrite = 1'b0;
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
        PerformanceCounterPlugin_logic_fsm_holdCsrWrite = 1'b0;
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_flusher_hits = {PerformanceCounterPlugin_logic_counters_instret_needFlush,PerformanceCounterPlugin_logic_counters_cycle_needFlush};
  assign PerformanceCounterPlugin_logic_flusher_hit = (|PerformanceCounterPlugin_logic_flusher_hits);
  assign PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input = PerformanceCounterPlugin_logic_flusher_hits;
  assign PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked = (PerformanceCounterPlugin_logic_flusher_hits_ohFirst_input & (~ _zz_PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked));
  assign PerformanceCounterPlugin_logic_flusher_oh = PerformanceCounterPlugin_logic_flusher_hits_ohFirst_masked;
  assign PerformanceCounterPlugin_logic_fsm_flusherCmd_valid = PerformanceCounterPlugin_logic_flusher_hit;
  assign PerformanceCounterPlugin_logic_fsm_flusherCmd_payload_oh = PerformanceCounterPlugin_logic_flusher_oh;
  assign PerformanceCounterPlugin_logic_csrDecode_addr = CsrAccessPlugin_bus_decode_address[1 : 0];
  always @(*) begin
    PerformanceCounterPlugin_logic_csrDecode_mok = 1'bx;
    case(PerformanceCounterPlugin_logic_csrDecode_addr)
      2'b00 : begin
        PerformanceCounterPlugin_logic_csrDecode_mok = PerformanceCounterPlugin_logic_counters_cycle_mcounteren;
      end
      2'b10 : begin
        PerformanceCounterPlugin_logic_csrDecode_mok = PerformanceCounterPlugin_logic_counters_instret_mcounteren;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    PerformanceCounterPlugin_logic_csrDecode_sok = 1'bx;
    case(PerformanceCounterPlugin_logic_csrDecode_addr)
      2'b00 : begin
        PerformanceCounterPlugin_logic_csrDecode_sok = PerformanceCounterPlugin_logic_counters_cycle_scounteren;
      end
      2'b10 : begin
        PerformanceCounterPlugin_logic_csrDecode_sok = PerformanceCounterPlugin_logic_counters_instret_scounteren;
      end
      default : begin
      end
    endcase
  end

  assign PerformanceCounterPlugin_logic_csrDecode_privOk = (&(PrivilegedPlugin_logic_harts_0_privilege | {PerformanceCounterPlugin_logic_csrDecode_mok,PerformanceCounterPlugin_logic_csrDecode_sok}));
  assign PerformanceCounterPlugin_logic_fsm_csrReadCmd_fire = (PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid && PerformanceCounterPlugin_logic_fsm_csrReadCmd_ready);
  assign PerformanceCounterPlugin_logic_csrRead_requested = (CsrAccessPlugin_bus_read_valid && REG_CSR_PerformanceCounterPlugin_logic_csrFilter);
  assign PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid = (PerformanceCounterPlugin_logic_csrRead_requested && (! PerformanceCounterPlugin_logic_csrRead_fired));
  assign PerformanceCounterPlugin_logic_fsm_csrReadCmd_payload_address = CsrAccessPlugin_bus_read_address[1 : 0];
  assign when_PerformanceCounterPlugin_l342 = ((! PerformanceCounterPlugin_logic_csrRead_fired) || (! PerformanceCounterPlugin_logic_fsm_done));
  assign PerformanceCounterPlugin_logic_fsm_csrWriteCmd_fire = (PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid && PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready);
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid = 1'b0;
    if(when_CsrAccessPlugin_l343_3) begin
      if(when_PerformanceCounterPlugin_l357) begin
        PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid = 1'b1;
      end
    end
  end

  assign PerformanceCounterPlugin_logic_fsm_csrWriteCmd_payload_address = CsrAccessPlugin_bus_write_address[1 : 0];
  assign CsrAccessPlugin_logic_fsm_wantExit = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_fsm_wantStart = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        CsrAccessPlugin_logic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign CsrAccessPlugin_logic_fsm_wantKill = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_fsm_interface_fire = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
        if(execute_ctrl2_down_isReady) begin
          CsrAccessPlugin_logic_fsm_interface_fire = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_logic_fsm_inject_csrAddress = execute_ctrl2_down_Decode_UOP_lane0[31 : 20];
  assign CsrAccessPlugin_logic_fsm_inject_immZero = (execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h0);
  assign CsrAccessPlugin_logic_fsm_inject_srcZero = (execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0 ? CsrAccessPlugin_logic_fsm_inject_immZero : (execute_ctrl2_down_Decode_UOP_lane0[19 : 15] == 5'h0));
  assign CsrAccessPlugin_logic_fsm_inject_csrWrite = (! (execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0 && CsrAccessPlugin_logic_fsm_inject_srcZero));
  assign CsrAccessPlugin_logic_fsm_inject_csrRead = (! ((! execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0) && (! execute_ctrl2_up_RD_ENABLE_lane0)));
  assign COMB_CSR_768 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h300);
  assign COMB_CSR_256 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h100);
  assign COMB_CSR_384 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h180);
  assign COMB_CSR_3008 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hbc0);
  assign COMB_CSR_1952 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a0);
  assign COMB_CSR_1953 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a1);
  assign COMB_CSR_1954 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h7a2);
  assign COMB_CSR_3857 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf11);
  assign COMB_CSR_3858 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf12);
  assign COMB_CSR_3859 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf13);
  assign COMB_CSR_3860 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hf14);
  assign COMB_CSR_769 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h301);
  assign COMB_CSR_834 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h342);
  assign COMB_CSR_836 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h344);
  assign COMB_CSR_772 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h304);
  assign COMB_CSR_770 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h302);
  assign COMB_CSR_771 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h303);
  assign COMB_CSR_322 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h142);
  assign COMB_CSR_260 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h104);
  assign COMB_CSR_324 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h144);
  assign COMB_CSR_3073 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc01);
  assign COMB_CSR_3201 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc81);
  assign COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h105),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h305)});
  assign COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h141),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h341)});
  assign COMB_CSR_774 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h306);
  assign COMB_CSR_262 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h106);
  assign COMB_CSR_800 = (CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h320);
  assign COMB_CSR_ = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h73f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc9f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb9f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h33f),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_),{_zz_COMB_CSR__1,{_zz_COMB_CSR__2,_zz_COMB_CSR__3}}}}}}});
  assign COMB_CSR_CsrRamPlugin_csrMapper_selFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc82),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb82),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc80),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb80),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc02),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb02),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter),{_zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_1,{_zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_2,_zz_COMB_CSR_CsrRamPlugin_csrMapper_selFilter_3}}}}}}}}});
  assign COMB_CSR_PerformanceCounterPlugin_logic_csrFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc82),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb82),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc80),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb80),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hc02),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'hb02),{(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter),(CsrAccessPlugin_logic_fsm_inject_csrAddress == _zz_COMB_CSR_PerformanceCounterPlugin_logic_csrFilter_1)}}}}}}});
  assign COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter = (|{(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h100),(CsrAccessPlugin_logic_fsm_inject_csrAddress == 12'h300)});
  assign CsrAccessPlugin_logic_fsm_inject_implemented = (|{COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter,{COMB_CSR_PerformanceCounterPlugin_logic_csrFilter,{COMB_CSR_CsrRamPlugin_csrMapper_selFilter,{COMB_CSR_,{COMB_CSR_800,{COMB_CSR_262,{COMB_CSR_774,{COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter,{COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter,{COMB_CSR_3201,{_zz_CsrAccessPlugin_logic_fsm_inject_implemented,_zz_CsrAccessPlugin_logic_fsm_inject_implemented_1}}}}}}}}}}});
  assign CsrAccessPlugin_logic_fsm_inject_onDecodeDo = ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_IDLE));
  assign when_CsrAccessPlugin_l155 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_384);
  assign when_MmuPlugin_l221 = (PrivilegedPlugin_logic_harts_0_m_status_tvm && (PrivilegedPlugin_logic_harts_0_privilege == 2'b01));
  assign when_CsrAccessPlugin_l155_1 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_3008);
  assign when_CsrAccessPlugin_l155_2 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_PerformanceCounterPlugin_logic_csrFilter);
  assign when_PerformanceCounterPlugin_l327 = (CsrAccessPlugin_bus_decode_address[9 : 8] == 2'b00);
  assign when_PerformanceCounterPlugin_l328 = (CsrAccessPlugin_bus_decode_write || (! PerformanceCounterPlugin_logic_csrDecode_privOk));
  assign when_CsrAccessPlugin_l155_3 = (CsrAccessPlugin_logic_fsm_inject_onDecodeDo && COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter);
  assign CsrAccessPlugin_logic_fsm_inject_trap = ((! CsrAccessPlugin_logic_fsm_inject_implemented) || CsrAccessPlugin_bus_decode_exception);
  assign CsrAccessPlugin_bus_decode_read = CsrAccessPlugin_logic_fsm_inject_csrRead;
  assign CsrAccessPlugin_bus_decode_write = CsrAccessPlugin_logic_fsm_inject_csrWrite;
  assign CsrAccessPlugin_bus_decode_address = CsrAccessPlugin_logic_fsm_inject_csrAddress;
  assign CsrAccessPlugin_logic_fsm_interface_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_rs1 = execute_ctrl2_up_integer_RS1_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_uop = execute_ctrl2_down_Decode_UOP_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_doImm = execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_doMask = execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_doClear = execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_rdEnable = execute_ctrl2_up_RD_ENABLE_lane0;
  assign CsrAccessPlugin_logic_fsm_interface_rdPhys = execute_ctrl2_down_RD_PHYS_lane0;
  assign CsrAccessPlugin_logic_fsm_inject_freeze = ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && (! CsrAccessPlugin_logic_fsm_inject_unfreeze));
  always @(*) begin
    CsrAccessPlugin_logic_flushPort_valid = 1'b0;
    if(CsrAccessPlugin_logic_fsm_inject_flushReg) begin
      CsrAccessPlugin_logic_flushPort_valid = 1'b1;
    end
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_flushPort_valid = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_flushPort_valid = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  assign CsrAccessPlugin_logic_flushPort_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign CsrAccessPlugin_logic_flushPort_payload_self = 1'b0;
  always @(*) begin
    CsrAccessPlugin_logic_trapPort_valid = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_trapPort_valid = 1'b1;
            end else begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_valid = 1'b1;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_trapPort_payload_exception = 1'b1;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_payload_exception = 1'b0;
              end
            end
          end
        end
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_trapPort_payload_code = 4'b0010;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              if(CsrAccessPlugin_logic_fsm_inject_busTrapReg) begin
                CsrAccessPlugin_logic_trapPort_payload_code = CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg;
              end
            end
          end
        end
      end
    endcase
  end

  assign CsrAccessPlugin_logic_trapPort_payload_tval = execute_ctrl2_down_Decode_UOP_lane0;
  assign CsrAccessPlugin_logic_trapPort_payload_arg = 3'b000;
  assign when_CsrAccessPlugin_l197 = (! execute_freeze_valid);
  always @(*) begin
    CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        CsrAccessPlugin_logic_fsm_readLogic_onReadsDo = CsrAccessPlugin_logic_fsm_interface_read;
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        if(when_CsrAccessPlugin_l296) begin
          CsrAccessPlugin_logic_fsm_readLogic_onReadsFireDo = CsrAccessPlugin_logic_fsm_interface_read;
        end
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_bus_read_valid = CsrAccessPlugin_logic_fsm_readLogic_onReadsDo;
  assign CsrAccessPlugin_bus_read_address = CsrAccessPlugin_logic_fsm_interface_uop[31 : 20];
  assign CsrAccessPlugin_bus_read_moving = (! CsrAccessPlugin_bus_read_halt);
  assign when_CsrAccessPlugin_l252 = (CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_CsrRamPlugin_csrMapper_selFilter);
  assign CsrAccessPlugin_logic_fsm_readLogic_csrValue = (((((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_20 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_31) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_40 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_47)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_54 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_64) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_74 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_85))) | (((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_96 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_107) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_118 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_127)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_138 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_149) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_160 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_171)))) | ((((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_180 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_184) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_186 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_188)) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_190 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_192) | (_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_194 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_196))) | ((_zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_198 | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_200) | _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_202)));
  assign CsrAccessPlugin_bus_read_data = CsrAccessPlugin_logic_fsm_readLogic_csrValue;
  always @(*) begin
    CsrAccessPlugin_bus_read_toWriteBits = CsrAccessPlugin_logic_fsm_readLogic_csrValue;
    if(when_CsrAccessPlugin_l279) begin
      if(when_CsrService_l198) begin
        CsrAccessPlugin_bus_read_toWriteBits[9 : 9] = PrivilegedPlugin_logic_harts_0_s_ip_seipSoft;
      end
    end
  end

  assign when_CsrAccessPlugin_l279 = (CsrAccessPlugin_logic_fsm_readLogic_onReadsDo && REG_CSR_836);
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue = REG_CSR_768;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_1 = REG_CSR_256;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_2 = REG_CSR_384;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_3 = REG_CSR_3008;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_6 = REG_CSR_836;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_8 = REG_CSR_772;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_11 = REG_CSR_771;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_17 = REG_CSR_774;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_18 = REG_CSR_262;
  assign _zz_CsrAccessPlugin_logic_fsm_readLogic_csrValue_19 = REG_CSR_800;
  assign when_CsrService_l198 = 1'b1;
  assign CsrAccessPlugin_bus_write_moving = (! CsrAccessPlugin_bus_write_halt);
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_mask = (CsrAccessPlugin_logic_fsm_interface_doImm ? _zz_CsrAccessPlugin_logic_fsm_writeLogic_alu_mask : CsrAccessPlugin_logic_fsm_interface_rs1);
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_masked = (CsrAccessPlugin_logic_fsm_interface_doClear ? (CsrAccessPlugin_logic_fsm_interface_aluInput & (~ CsrAccessPlugin_logic_fsm_writeLogic_alu_mask)) : (CsrAccessPlugin_logic_fsm_interface_aluInput | CsrAccessPlugin_logic_fsm_writeLogic_alu_mask));
  assign CsrAccessPlugin_logic_fsm_writeLogic_alu_result = (CsrAccessPlugin_logic_fsm_interface_doMask ? CsrAccessPlugin_logic_fsm_writeLogic_alu_masked : CsrAccessPlugin_logic_fsm_writeLogic_alu_mask);
  always @(*) begin
    CsrAccessPlugin_bus_write_bits = CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
    if(when_CsrAccessPlugin_l343) begin
      CsrAccessPlugin_bus_write_bits[1 : 0] = 2'b00;
    end
    if(when_CsrAccessPlugin_l343_1) begin
      CsrAccessPlugin_bus_write_bits[1 : 0] = 2'b00;
    end
  end

  assign CsrAccessPlugin_bus_write_address = CsrAccessPlugin_logic_fsm_interface_uop[31 : 20];
  always @(*) begin
    CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
        CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo = CsrAccessPlugin_logic_fsm_interface_write;
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = 1'b0;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
        if(when_CsrAccessPlugin_l325) begin
          CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo = CsrAccessPlugin_logic_fsm_interface_write;
        end
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrAccessPlugin_bus_write_valid = CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo;
  assign when_CsrService_l176 = 1'b1;
  assign when_CsrAccessPlugin_l346 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_768);
  assign switch_PrivilegedPlugin_l549 = CsrAccessPlugin_bus_write_bits[12 : 11];
  assign when_CsrAccessPlugin_l346_1 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_256);
  assign when_CsrAccessPlugin_l353 = ((|((MmuPlugin_logic_satpModeWrite != 1'b0) && (MmuPlugin_logic_satpModeWrite != 1'b1))) == 1'b0);
  assign when_CsrAccessPlugin_l346_2 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_384);
  assign when_CsrAccessPlugin_l346_3 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_3008);
  assign when_CsrAccessPlugin_l346_4 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_834);
  assign when_CsrAccessPlugin_l346_5 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_836);
  assign when_CsrAccessPlugin_l346_6 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_772);
  assign when_CsrAccessPlugin_l346_7 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_770);
  assign when_CsrAccessPlugin_l346_8 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_771);
  assign when_CsrAccessPlugin_l346_9 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_322);
  assign when_CsrAccessPlugin_l346_10 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_260);
  assign when_CsrAccessPlugin_l346_11 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_324);
  assign when_CsrAccessPlugin_l343 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter);
  assign when_CsrAccessPlugin_l343_1 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter);
  assign when_CsrAccessPlugin_l346_12 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_774);
  assign when_CsrAccessPlugin_l346_13 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_262);
  assign when_CsrAccessPlugin_l346_14 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesFireDo && REG_CSR_800);
  assign when_CsrAccessPlugin_l343_2 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_CsrRamPlugin_csrMapper_selFilter);
  assign when_CsrAccessPlugin_l343_3 = (CsrAccessPlugin_logic_fsm_writeLogic_onWritesDo && REG_CSR_PerformanceCounterPlugin_logic_csrFilter);
  assign when_PerformanceCounterPlugin_l357 = (! PerformanceCounterPlugin_logic_csrWrite_fired);
  assign when_PerformanceCounterPlugin_l359 = (! PerformanceCounterPlugin_logic_fsm_csrWriteCmd_ready);
  assign CsrAccessPlugin_logic_wbWi_valid = execute_ctrl3_down_CsrAccessPlugin_SEL_lane0;
  assign CsrAccessPlugin_logic_wbWi_payload = CsrAccessPlugin_logic_fsm_interface_csrValue;
  assign FetchL1Plugin_pmaBuilder_addressBits = FetchL1Plugin_logic_ctrl_pmaPort_cmd_address;
  assign _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io = ((FetchL1Plugin_pmaBuilder_addressBits & 32'h0) == 32'h0);
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit = _zz_FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit[0];
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit = (|1'b1);
  assign FetchL1Plugin_pmaBuilder_onTransfers_0_hit = (FetchL1Plugin_pmaBuilder_onTransfers_0_argsHit && FetchL1Plugin_pmaBuilder_onTransfers_0_addressHit);
  assign FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault = (! ((|{((FetchL1Plugin_pmaBuilder_addressBits & 32'hf0000000) == 32'h40000000),{((FetchL1Plugin_pmaBuilder_addressBits & 32'hffff0000) == 32'h0),{((FetchL1Plugin_pmaBuilder_addressBits & _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault) == 32'h10000000),((FetchL1Plugin_pmaBuilder_addressBits & _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_fault_1) == 32'h10001000)}}}) && (|FetchL1Plugin_pmaBuilder_onTransfers_0_hit)));
  assign FetchL1Plugin_logic_ctrl_pmaPort_rsp_io = (! _zz_FetchL1Plugin_logic_ctrl_pmaPort_rsp_io_1[0]);
  assign LsuPlugin_pmaBuilder_l1_addressBits = LsuPlugin_logic_onPma_cached_cmd_address;
  assign LsuPlugin_pmaBuilder_l1_argsBits = LsuPlugin_logic_onPma_cached_cmd_op;
  assign _zz_LsuPlugin_logic_onPma_cached_rsp_io = ((LsuPlugin_pmaBuilder_l1_addressBits & 32'h0) == 32'h0);
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit = _zz_LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit[0];
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit = (|((LsuPlugin_pmaBuilder_l1_argsBits & 1'b0) == 1'b0));
  assign LsuPlugin_pmaBuilder_l1_onTransfers_0_hit = (LsuPlugin_pmaBuilder_l1_onTransfers_0_argsHit && LsuPlugin_pmaBuilder_l1_onTransfers_0_addressHit);
  assign LsuPlugin_logic_onPma_cached_rsp_fault = (! ((|{((LsuPlugin_pmaBuilder_l1_addressBits & 32'hf0000000) == 32'h40000000),{((LsuPlugin_pmaBuilder_l1_addressBits & 32'hff000000) == 32'h01000000),{((LsuPlugin_pmaBuilder_l1_addressBits & _zz_LsuPlugin_logic_onPma_cached_rsp_fault) == 32'h0),{(_zz_LsuPlugin_logic_onPma_cached_rsp_fault_1 == _zz_LsuPlugin_logic_onPma_cached_rsp_fault_2),(_zz_LsuPlugin_logic_onPma_cached_rsp_fault_3 == _zz_LsuPlugin_logic_onPma_cached_rsp_fault_4)}}}}) && (|LsuPlugin_pmaBuilder_l1_onTransfers_0_hit)));
  assign LsuPlugin_logic_onPma_cached_rsp_io = (! _zz_LsuPlugin_logic_onPma_cached_rsp_io_1[0]);
  assign LsuPlugin_pmaBuilder_io_addressBits = LsuPlugin_logic_onPma_io_cmd_address;
  assign LsuPlugin_pmaBuilder_io_argsBits = {LsuPlugin_logic_onPma_io_cmd_size,LsuPlugin_logic_onPma_io_cmd_op};
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit = _zz_LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit[0];
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit = (|{((LsuPlugin_pmaBuilder_io_argsBits & 3'b100) == 3'b100),((LsuPlugin_pmaBuilder_io_argsBits & 3'b001) == 3'b000)});
  assign LsuPlugin_pmaBuilder_io_onTransfers_0_hit = (LsuPlugin_pmaBuilder_io_onTransfers_0_argsHit && LsuPlugin_pmaBuilder_io_onTransfers_0_addressHit);
  assign _zz_LsuPlugin_logic_onPma_io_rsp_io = ((LsuPlugin_pmaBuilder_io_addressBits & 32'h80000000) == 32'h0);
  assign LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit = _zz_LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit[0];
  assign LsuPlugin_pmaBuilder_io_onTransfers_1_argsHit = (|((LsuPlugin_pmaBuilder_io_argsBits & 3'b000) == 3'b000));
  assign LsuPlugin_pmaBuilder_io_onTransfers_1_hit = (LsuPlugin_pmaBuilder_io_onTransfers_1_argsHit && LsuPlugin_pmaBuilder_io_onTransfers_1_addressHit);
  assign LsuPlugin_logic_onPma_io_rsp_fault = (! ((|{((LsuPlugin_pmaBuilder_io_addressBits & 32'hff000000) == 32'h01000000),{((LsuPlugin_pmaBuilder_io_addressBits & _zz_LsuPlugin_logic_onPma_io_rsp_fault) == 32'hf0c00000),{(_zz_LsuPlugin_logic_onPma_io_rsp_fault_1 == _zz_LsuPlugin_logic_onPma_io_rsp_fault_2),{_zz_LsuPlugin_logic_onPma_io_rsp_fault_3,{_zz_LsuPlugin_logic_onPma_io_rsp_fault_4,_zz_LsuPlugin_logic_onPma_io_rsp_fault_5}}}}}) && (|{LsuPlugin_pmaBuilder_io_onTransfers_1_hit,LsuPlugin_pmaBuilder_io_onTransfers_0_hit})));
  assign LsuPlugin_logic_onPma_io_rsp_io = (! _zz_LsuPlugin_logic_onPma_io_rsp_io_1[0]);
  assign CsrRamPlugin_logic_writeLogic_hits = {CsrRamPlugin_setup_initPort_valid,{CsrRamPlugin_csrMapper_write_valid,{TrapPlugin_logic_harts_0_crsPorts_write_valid,PerformanceCounterPlugin_logic_writePort_valid}}};
  assign CsrRamPlugin_logic_writeLogic_hit = (|CsrRamPlugin_logic_writeLogic_hits);
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_input = CsrRamPlugin_logic_writeLogic_hits;
  assign CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_writeLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_writeLogic_oh = CsrRamPlugin_logic_writeLogic_hits_ohFirst_masked;
  assign _zz_PerformanceCounterPlugin_logic_writePort_ready = CsrRamPlugin_logic_writeLogic_oh[0];
  assign _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready = CsrRamPlugin_logic_writeLogic_oh[1];
  assign _zz_CsrRamPlugin_csrMapper_write_ready = CsrRamPlugin_logic_writeLogic_oh[2];
  assign _zz_CsrRamPlugin_setup_initPort_ready = CsrRamPlugin_logic_writeLogic_oh[3];
  assign CsrRamPlugin_logic_writeLogic_port_valid = CsrRamPlugin_logic_writeLogic_hit;
  assign CsrRamPlugin_logic_writeLogic_port_payload_address = (((_zz_PerformanceCounterPlugin_logic_writePort_ready ? PerformanceCounterPlugin_logic_writePort_address : 4'b0000) | (_zz_TrapPlugin_logic_harts_0_crsPorts_write_ready ? TrapPlugin_logic_harts_0_crsPorts_write_address : 4'b0000)) | ((_zz_CsrRamPlugin_csrMapper_write_ready ? CsrRamPlugin_csrMapper_write_address : 4'b0000) | (_zz_CsrRamPlugin_setup_initPort_ready ? CsrRamPlugin_setup_initPort_address : 4'b0000)));
  assign CsrRamPlugin_logic_writeLogic_port_payload_data = (((_zz_PerformanceCounterPlugin_logic_writePort_ready ? PerformanceCounterPlugin_logic_writePort_data : 32'h0) | (_zz_TrapPlugin_logic_harts_0_crsPorts_write_ready ? TrapPlugin_logic_harts_0_crsPorts_write_data : 32'h0)) | ((_zz_CsrRamPlugin_csrMapper_write_ready ? CsrRamPlugin_csrMapper_write_data : 32'h0) | (_zz_CsrRamPlugin_setup_initPort_ready ? CsrRamPlugin_setup_initPort_data : 32'h0)));
  assign PerformanceCounterPlugin_logic_writePort_ready = _zz_PerformanceCounterPlugin_logic_writePort_ready;
  assign TrapPlugin_logic_harts_0_crsPorts_write_ready = _zz_TrapPlugin_logic_harts_0_crsPorts_write_ready;
  assign CsrRamPlugin_csrMapper_write_ready = _zz_CsrRamPlugin_csrMapper_write_ready;
  assign CsrRamPlugin_setup_initPort_ready = _zz_CsrRamPlugin_setup_initPort_ready;
  assign CsrRamPlugin_logic_readLogic_hits = {CsrRamPlugin_csrMapper_read_valid,{TrapPlugin_logic_harts_0_crsPorts_read_valid,PerformanceCounterPlugin_logic_readPort_valid}};
  assign CsrRamPlugin_logic_readLogic_hit = (|CsrRamPlugin_logic_readLogic_hits);
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_input = CsrRamPlugin_logic_readLogic_hits;
  assign CsrRamPlugin_logic_readLogic_hits_ohFirst_masked = (CsrRamPlugin_logic_readLogic_hits_ohFirst_input & (~ _zz_CsrRamPlugin_logic_readLogic_hits_ohFirst_masked));
  assign CsrRamPlugin_logic_readLogic_oh = CsrRamPlugin_logic_readLogic_hits_ohFirst_masked;
  assign _zz_CsrRamPlugin_logic_readLogic_sel = CsrRamPlugin_logic_readLogic_oh[1];
  assign _zz_CsrRamPlugin_logic_readLogic_sel_1 = CsrRamPlugin_logic_readLogic_oh[2];
  assign CsrRamPlugin_logic_readLogic_sel = {_zz_CsrRamPlugin_logic_readLogic_sel_1,_zz_CsrRamPlugin_logic_readLogic_sel};
  assign CsrRamPlugin_logic_readLogic_port_rsp = CsrRamPlugin_logic_mem_spinal_port1;
  assign CsrRamPlugin_logic_readLogic_port_cmd_valid = (((|CsrRamPlugin_logic_readLogic_oh) && (! CsrRamPlugin_logic_writeLogic_port_valid)) && (! CsrRamPlugin_logic_readLogic_busy));
  assign CsrRamPlugin_logic_readLogic_port_cmd_payload = _zz_CsrRamPlugin_logic_readLogic_port_cmd_payload;
  assign PerformanceCounterPlugin_logic_readPort_ready = CsrRamPlugin_logic_readLogic_ohReg[0];
  assign TrapPlugin_logic_harts_0_crsPorts_read_ready = CsrRamPlugin_logic_readLogic_ohReg[1];
  assign CsrRamPlugin_csrMapper_read_ready = CsrRamPlugin_logic_readLogic_ohReg[2];
  assign PerformanceCounterPlugin_logic_readPort_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign TrapPlugin_logic_harts_0_crsPorts_read_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign CsrRamPlugin_csrMapper_read_data = CsrRamPlugin_logic_readLogic_port_rsp;
  assign CsrRamPlugin_logic_flush_done = CsrRamPlugin_logic_flush_counter[4];
  assign CsrRamPlugin_setup_initPort_valid = (! CsrRamPlugin_logic_flush_done);
  assign CsrRamPlugin_setup_initPort_address = CsrRamPlugin_logic_flush_counter[3:0];
  assign CsrRamPlugin_setup_initPort_data = 32'h0;
  assign execute_lane0_bypasser_integer_RS1_port_valid = (! execute_freeze_valid);
  assign execute_lane0_bypasser_integer_RS1_port_address = execute_ctrl0_down_RS1_PHYS_lane0;
  always @(*) begin
    execute_lane0_bypasser_integer_RS1_bypassEnables[0] = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS1_bypassEnables[1] = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS1_bypassEnables[2] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS1_bypassEnables[3] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS1_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS1_bypassEnables[4] = 1'b1;
  end

  assign _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 = execute_lane0_bypasser_integer_RS1_bypassEnables;
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[0];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[1];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[2];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[3];
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 = _zz_execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0[4];
  always @(*) begin
    _zz_execute_lane0_bypasser_integer_RS1_sel[0] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane0_bypasser_integer_RS1_sel[1] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0));
    _zz_execute_lane0_bypasser_integer_RS1_sel[2] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1));
    _zz_execute_lane0_bypasser_integer_RS1_sel[3] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2));
    _zz_execute_lane0_bypasser_integer_RS1_sel[4] = (execute_lane0_bypasser_integer_RS1_bypassEnables_bools_4 && (! execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3));
  end

  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_1 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0});
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_2 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0}});
  assign execute_lane0_bypasser_integer_RS1_bypassEnables_range_0_to_3 = (|{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_3,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS1_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS1_bypassEnables_bools_0}}});
  assign execute_lane0_bypasser_integer_RS1_sel = _zz_execute_lane0_bypasser_integer_RS1_sel;
  assign _zz_execute_ctrl1_down_integer_RS1_lane0 = execute_lane0_bypasser_integer_RS1_sel[4 : 1];
  always @(*) begin
    _zz_execute_ctrl1_down_integer_RS1_lane0_1 = (((_zz_execute_ctrl1_down_integer_RS1_lane0[0] ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_execute_ctrl1_down_integer_RS1_lane0[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_execute_ctrl1_down_integer_RS1_lane0[2] ? execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_execute_ctrl1_down_integer_RS1_lane0[3] ? execute_lane0_bypasser_integer_RS1_port_data : 32'h0)));
    if(when_ExecuteLanePlugin_l196) begin
      _zz_execute_ctrl1_down_integer_RS1_lane0_1 = execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign execute_ctrl1_down_integer_RS1_lane0 = _zz_execute_ctrl1_down_integer_RS1_lane0_1;
  assign when_ExecuteLanePlugin_l196 = execute_lane0_bypasser_integer_RS1_sel[0];
  assign execute_lane0_bypasser_integer_RS2_port_valid = (! execute_freeze_valid);
  assign execute_lane0_bypasser_integer_RS2_port_address = execute_ctrl0_down_RS2_PHYS_lane0;
  always @(*) begin
    execute_lane0_bypasser_integer_RS2_bypassEnables[0] = (((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_up_RD_ENABLE_lane0) && (execute_ctrl2_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS2_bypassEnables[1] = (((execute_ctrl3_up_LANE_SEL_lane0 && execute_ctrl3_up_RD_ENABLE_lane0) && (execute_ctrl3_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS2_bypassEnables[2] = (((execute_ctrl4_up_LANE_SEL_lane0 && execute_ctrl4_up_RD_ENABLE_lane0) && (execute_ctrl4_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS2_bypassEnables[3] = (((execute_ctrl5_up_LANE_SEL_lane0 && execute_ctrl5_up_RD_ENABLE_lane0) && (execute_ctrl5_down_RD_PHYS_lane0 == execute_ctrl1_down_RS2_PHYS_lane0)) && 1'b1);
    execute_lane0_bypasser_integer_RS2_bypassEnables[4] = 1'b1;
  end

  assign _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 = execute_lane0_bypasser_integer_RS2_bypassEnables;
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[0];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[1];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[2];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[3];
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 = _zz_execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0[4];
  always @(*) begin
    _zz_execute_lane0_bypasser_integer_RS2_sel[0] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0 && (! 1'b0));
    _zz_execute_lane0_bypasser_integer_RS2_sel[1] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0));
    _zz_execute_lane0_bypasser_integer_RS2_sel[2] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1));
    _zz_execute_lane0_bypasser_integer_RS2_sel[3] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2));
    _zz_execute_lane0_bypasser_integer_RS2_sel[4] = (execute_lane0_bypasser_integer_RS2_bypassEnables_bools_4 && (! execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3));
  end

  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_1 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0});
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_2 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0}});
  assign execute_lane0_bypasser_integer_RS2_bypassEnables_range_0_to_3 = (|{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_3,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_2,{execute_lane0_bypasser_integer_RS2_bypassEnables_bools_1,execute_lane0_bypasser_integer_RS2_bypassEnables_bools_0}}});
  assign execute_lane0_bypasser_integer_RS2_sel = _zz_execute_lane0_bypasser_integer_RS2_sel;
  assign _zz_execute_ctrl1_down_integer_RS2_lane0 = execute_lane0_bypasser_integer_RS2_sel[4 : 1];
  always @(*) begin
    _zz_execute_ctrl1_down_integer_RS2_lane0_1 = (((_zz_execute_ctrl1_down_integer_RS2_lane0[0] ? execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_execute_ctrl1_down_integer_RS2_lane0[1] ? execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0)) | ((_zz_execute_ctrl1_down_integer_RS2_lane0[2] ? execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 : 32'h0) | (_zz_execute_ctrl1_down_integer_RS2_lane0[3] ? execute_lane0_bypasser_integer_RS2_port_data : 32'h0)));
    if(when_ExecuteLanePlugin_l196_1) begin
      _zz_execute_ctrl1_down_integer_RS2_lane0_1 = execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
  end

  assign execute_ctrl1_down_integer_RS2_lane0 = _zz_execute_ctrl1_down_integer_RS2_lane0_1;
  assign when_ExecuteLanePlugin_l196_1 = execute_lane0_bypasser_integer_RS2_sel[0];
  assign execute_lane0_logic_completions_onCtrl_0_port_valid = (((execute_ctrl2_down_LANE_SEL_lane0 && execute_ctrl2_down_isReady) && (! execute_lane0_ctrls_2_downIsCancel)) && execute_ctrl2_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_uopId = execute_ctrl2_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_trap = execute_ctrl2_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_0_port_payload_commit = execute_ctrl2_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_valid = (((execute_ctrl3_down_LANE_SEL_lane0 && execute_ctrl3_down_isReady) && (! execute_lane0_ctrls_3_downIsCancel)) && execute_ctrl3_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_uopId = execute_ctrl3_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_trap = execute_ctrl3_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_1_port_payload_commit = execute_ctrl3_down_COMMIT_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_valid = (((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0);
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_trap = execute_ctrl4_down_TRAP_lane0;
  assign execute_lane0_logic_completions_onCtrl_2_port_payload_commit = execute_ctrl4_down_COMMIT_lane0;
  assign execute_lane0_logic_decoding_decodingBits = execute_ctrl1_down_Decode_UOP_lane0;
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h0000004c) == 32'h00000004);
  always @(*) begin
    execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000050) == 32'h00000040);
  always @(*) begin
    execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_BranchPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_BranchPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_MulPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_MulPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_DivPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_DivPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_early0_EnvPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h0000000c) == 32'h00000008);
  always @(*) begin
    execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0 = _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_SEL_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_CsrAccessPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_AguPlugin_SEL_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000058) == 32'h0);
  always @(*) begin
    execute_ctrl1_down_AguPlugin_SEL_lane0 = _zz_execute_ctrl1_down_AguPlugin_SEL_lane0_1[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_AguPlugin_SEL_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000028) == 32'h0);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h0000000c) == 32'h00000004);
  assign _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00002008) == 32'h00002008);
  always @(*) begin
    execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = _zz_execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0_1[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 32'h02003010) == 32'h00000010);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 32'h10003010) == 32'h10000010);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 32'h02000050) == 32'h00000010);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_4 = ((execute_lane0_logic_decoding_decodingBits & 32'h00001044) == 32'h00001004);
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000030) == 32'h00000010);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_2_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_2_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_2_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 32'h0200402c) == 32'h02004020);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 32'h00001040) == 32'h00001040);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_3 = ((execute_lane0_logic_decoding_decodingBits & 32'h00002040) == 32'h00002040);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_3_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_3_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_3_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h02004064) == 32'h02000020);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_1 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000054) == 32'h0);
  assign _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 32'h00001050) == 32'h0);
  always @(*) begin
    execute_ctrl1_down_COMPLETION_AT_4_lane0 = _zz_execute_ctrl1_down_COMPLETION_AT_4_lane0[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_COMPLETION_AT_4_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0_5[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0_4[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = 1'b0;
    end
  end

  always @(*) begin
    execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = _zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0_3[0];
    if(execute_ctrl1_down_TRAP_lane0) begin
      execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = 1'b0;
    end
  end

  assign _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00006000) == 32'h0);
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000004) == 32'h00000004);
  assign execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0_1[0];
  assign execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0[0];
  assign _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00004000) == 32'h0);
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00001000) == 32'h00001000);
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1 = {(|{_zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0,{_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0,_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0}}),(|{_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0,{_zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h00003000) == 32'h00002000)}})};
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_1;
  assign _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = _zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0_2;
  assign _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_2 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000040) == 32'h00000040);
  assign execute_ctrl1_down_SrcStageables_REVERT_lane0 = _zz_execute_ctrl1_down_SrcStageables_REVERT_lane0[0];
  assign execute_ctrl1_down_SrcStageables_ZERO_lane0 = _zz_execute_ctrl1_down_SrcStageables_ZERO_lane0[0];
  assign execute_ctrl1_down_early0_SrcPlugin_logic_SRC1_CTRL_lane0 = (|_zz_execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0);
  assign execute_ctrl1_down_early0_SrcPlugin_logic_SRC2_CTRL_lane0 = {(|{_zz_execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0,((execute_lane0_logic_decoding_decodingBits & 32'h00000070) == 32'h00000020)}),(|{((execute_lane0_logic_decoding_decodingBits & 32'h00000050) == 32'h0),((execute_lane0_logic_decoding_decodingBits & 32'h00000024) == 32'h0)})};
  assign execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0[0];
  assign _zz_execute_ctrl1_down_AguPlugin_STORE_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h10000020) == 32'h00000020);
  assign execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = {(|{((execute_lane0_logic_decoding_decodingBits & 32'h00000010) == 32'h00000010),{((execute_lane0_logic_decoding_decodingBits & _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0) == 32'h00002000),{_zz_execute_ctrl1_down_AguPlugin_STORE_lane0,(_zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_1 == _zz_execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0_2)}}}),(|((execute_lane0_logic_decoding_decodingBits & 32'h00001010) == 32'h00001000))};
  assign execute_ctrl1_down_BYPASSED_AT_2_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_2_lane0[0];
  assign execute_ctrl1_down_BYPASSED_AT_3_lane0 = _zz_execute_ctrl1_down_BYPASSED_AT_3_lane0_3[0];
  assign execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0[0];
  assign execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0 = _zz_execute_ctrl1_down_MAY_FLUSH_PRECISE_4_lane0[0];
  assign execute_ctrl1_down_SrcStageables_UNSIGNED_lane0 = _zz_execute_ctrl1_down_SrcStageables_UNSIGNED_lane0[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0_1[0];
  assign execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0 = _zz_execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0[0];
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1 = {(|_zz_execute_ctrl1_down_BYPASSED_AT_3_lane0),(|((execute_lane0_logic_decoding_decodingBits & 32'h00000008) == 32'h00000008))};
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_1;
  assign _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
  assign execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0 = _zz_execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0_2;
  assign execute_ctrl1_down_CfuPlugin_logic_CFU_ENCODING_lane0 = (|((execute_lane0_logic_decoding_decodingBits & 32'h0) == 32'h0));
  assign _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_1 = (|((execute_lane0_logic_decoding_decodingBits & 32'h00000020) == 32'h00000020));
  assign _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0 = _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_1;
  assign _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_2 = _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0;
  assign execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0 = _zz_execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0_2;
  assign _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00002000) == 32'h00002000);
  assign execute_ctrl1_down_MulPlugin_HIGH_lane0 = _zz_execute_ctrl1_down_MulPlugin_HIGH_lane0[0];
  assign execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0[0];
  assign execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = _zz_execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0_1[0];
  assign execute_ctrl1_down_DivPlugin_REM_lane0 = _zz_execute_ctrl1_down_DivPlugin_REM_lane0[0];
  assign execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0[0];
  assign execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0_1[0];
  assign execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0 = _zz_execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_LOAD_lane0 = _zz_execute_ctrl1_down_AguPlugin_LOAD_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_STORE_lane0 = _zz_execute_ctrl1_down_AguPlugin_STORE_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_ATOMIC_lane0 = _zz_execute_ctrl1_down_AguPlugin_ATOMIC_lane0_1[0];
  assign execute_ctrl1_down_AguPlugin_FLOAT_lane0 = _zz_execute_ctrl1_down_AguPlugin_FLOAT_lane0[0];
  assign execute_ctrl1_down_AguPlugin_CLEAN_lane0 = _zz_execute_ctrl1_down_AguPlugin_CLEAN_lane0[0];
  assign execute_ctrl1_down_AguPlugin_INVALIDATE_lane0 = _zz_execute_ctrl1_down_AguPlugin_INVALIDATE_lane0[0];
  assign execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = _zz_execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0[0];
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0 = ((execute_lane0_logic_decoding_decodingBits & 32'h00000040) == 32'h0);
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2 = {(|{((execute_lane0_logic_decoding_decodingBits & _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2) == 32'h02000000),((execute_lane0_logic_decoding_decodingBits & _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_1) == 32'h10000000)}),{(|{_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0,(_zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_2 == _zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_3)}),(|{_zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0,{_zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_4,_zz__zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2_5}})}};
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1 = _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_2;
  assign _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3 = _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_1;
  assign execute_ctrl1_down_early0_EnvPlugin_OP_lane0 = _zz_execute_ctrl1_down_early0_EnvPlugin_OP_lane0_3;
  assign when_ExecuteLanePlugin_l306 = (|{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}});
  assign execute_lane0_ctrls_0_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_0_upIsCancel = when_ExecuteLanePlugin_l306;
  assign when_ExecuteLanePlugin_l306_1 = (|{(early0_EnvPlugin_logic_flushPort_valid && 1'b1),{(CsrAccessPlugin_logic_flushPort_valid && 1'b1),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}});
  assign execute_lane0_ctrls_1_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_1_upIsCancel = when_ExecuteLanePlugin_l306_1;
  assign when_ExecuteLanePlugin_l306_2 = (|{((early0_EnvPlugin_logic_flushPort_valid && 1'b1) && (1'b0 || (1'b1 && early0_EnvPlugin_logic_flushPort_payload_self))),{((CsrAccessPlugin_logic_flushPort_valid && 1'b1) && (1'b0 || (_zz_when_ExecuteLanePlugin_l306_2 && CsrAccessPlugin_logic_flushPort_payload_self))),{(early0_BranchPlugin_logic_flushPort_valid && 1'b1),(LsuPlugin_logic_flushPort_valid && 1'b1)}}});
  assign execute_lane0_ctrls_2_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_2_upIsCancel = when_ExecuteLanePlugin_l306_2;
  assign when_ExecuteLanePlugin_l306_3 = (|{((early0_BranchPlugin_logic_flushPort_valid && 1'b1) && (1'b0 || (1'b1 && early0_BranchPlugin_logic_flushPort_payload_self))),(LsuPlugin_logic_flushPort_valid && 1'b1)});
  assign execute_lane0_ctrls_3_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_3_upIsCancel = when_ExecuteLanePlugin_l306_3;
  assign when_ExecuteLanePlugin_l306_4 = (|((LsuPlugin_logic_flushPort_valid && 1'b1) && (1'b0 || (1'b1 && LsuPlugin_logic_flushPort_payload_self))));
  assign execute_lane0_ctrls_4_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_4_upIsCancel = when_ExecuteLanePlugin_l306_4;
  assign execute_lane0_ctrls_5_downIsCancel = 1'b0;
  assign execute_lane0_ctrls_5_upIsCancel = 1'b0;
  assign execute_lane0_logic_trapPending[0] = (|{((execute_ctrl4_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl4_down_TRAP_lane0),{((execute_ctrl3_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl3_down_TRAP_lane0),{((execute_ctrl2_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl2_down_TRAP_lane0),((execute_ctrl1_up_LANE_SEL_lane0 && 1'b1) && execute_ctrl1_down_TRAP_lane0)}}});
  assign execute_ctrl2_up_COMMIT_lane0 = (! execute_ctrl2_up_TRAP_lane0);
  assign WhiteboxerPlugin_logic_csr_access_valid = CsrAccessPlugin_logic_fsm_interface_fire;
  assign WhiteboxerPlugin_logic_csr_access_payload_uopId = CsrAccessPlugin_logic_fsm_interface_uopId;
  assign WhiteboxerPlugin_logic_csr_access_payload_address = _zz_WhiteboxerPlugin_logic_csr_access_payload_address[31 : 20];
  assign WhiteboxerPlugin_logic_csr_access_payload_write = CsrAccessPlugin_logic_fsm_interface_onWriteBits;
  assign WhiteboxerPlugin_logic_csr_access_payload_read = CsrAccessPlugin_logic_fsm_interface_csrValue;
  assign WhiteboxerPlugin_logic_csr_access_payload_writeDone = CsrAccessPlugin_logic_fsm_interface_write;
  assign WhiteboxerPlugin_logic_csr_access_payload_readDone = CsrAccessPlugin_logic_fsm_interface_read;
  assign WhiteboxerPlugin_logic_csr_port_valid = WhiteboxerPlugin_logic_csr_access_valid;
  assign WhiteboxerPlugin_logic_csr_port_payload_uopId = WhiteboxerPlugin_logic_csr_access_payload_uopId;
  assign WhiteboxerPlugin_logic_csr_port_payload_address = WhiteboxerPlugin_logic_csr_access_payload_address;
  assign WhiteboxerPlugin_logic_csr_port_payload_write = WhiteboxerPlugin_logic_csr_access_payload_write;
  assign WhiteboxerPlugin_logic_csr_port_payload_read = WhiteboxerPlugin_logic_csr_access_payload_read;
  assign WhiteboxerPlugin_logic_csr_port_payload_writeDone = WhiteboxerPlugin_logic_csr_access_payload_writeDone;
  assign WhiteboxerPlugin_logic_csr_port_payload_readDone = WhiteboxerPlugin_logic_csr_access_payload_readDone;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_valid = lane0_integer_WriteBackPlugin_logic_stages_0_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_0_payload_data = lane0_integer_WriteBackPlugin_logic_stages_0_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_valid = lane0_integer_WriteBackPlugin_logic_stages_1_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_1_payload_data = lane0_integer_WriteBackPlugin_logic_stages_1_write_payload_data;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_valid = lane0_integer_WriteBackPlugin_logic_stages_2_write_valid;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_payload_uopId = lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_uopId;
  assign WhiteboxerPlugin_logic_rfWrites_ports_2_payload_data = lane0_integer_WriteBackPlugin_logic_stages_2_write_payload_data;
  assign WhiteboxerPlugin_logic_completions_ports_0_valid = DecoderPlugin_logic_laneLogic_0_completionPort_valid;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_uopId = DecoderPlugin_logic_laneLogic_0_completionPort_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_trap = DecoderPlugin_logic_laneLogic_0_completionPort_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_0_payload_commit = DecoderPlugin_logic_laneLogic_0_completionPort_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_1_valid = execute_lane0_logic_completions_onCtrl_0_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_uopId = execute_lane0_logic_completions_onCtrl_0_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_trap = execute_lane0_logic_completions_onCtrl_0_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_1_payload_commit = execute_lane0_logic_completions_onCtrl_0_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_2_valid = execute_lane0_logic_completions_onCtrl_1_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_uopId = execute_lane0_logic_completions_onCtrl_1_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_trap = execute_lane0_logic_completions_onCtrl_1_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_2_payload_commit = execute_lane0_logic_completions_onCtrl_1_port_payload_commit;
  assign WhiteboxerPlugin_logic_completions_ports_3_valid = execute_lane0_logic_completions_onCtrl_2_port_valid;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_uopId = execute_lane0_logic_completions_onCtrl_2_port_payload_uopId;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_trap = execute_lane0_logic_completions_onCtrl_2_port_payload_trap;
  assign WhiteboxerPlugin_logic_completions_ports_3_payload_commit = execute_lane0_logic_completions_onCtrl_2_port_payload_commit;
  assign WhiteboxerPlugin_logic_commits_ports_0_oh_0 = ((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_COMMIT_lane0) && 1'b1);
  assign WhiteboxerPlugin_logic_commits_ports_0_valid = (|WhiteboxerPlugin_logic_commits_ports_0_oh_0);
  assign WhiteboxerPlugin_logic_commits_ports_0_pc = (WhiteboxerPlugin_logic_commits_ports_0_oh_0 ? execute_ctrl4_down_PC_lane0 : 32'h0);
  assign WhiteboxerPlugin_logic_commits_ports_0_uop = (WhiteboxerPlugin_logic_commits_ports_0_oh_0 ? execute_ctrl4_down_Decode_UOP_lane0 : 32'h0);
  assign WhiteboxerPlugin_logic_reschedules_flushes_0_valid = BtbPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_0_payload_self = BtbPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_valid = LsuPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_uopId = LsuPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_1_payload_self = LsuPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_valid = early0_BranchPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_uopId = early0_BranchPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_2_payload_self = early0_BranchPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_valid = CsrAccessPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_uopId = CsrAccessPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_3_payload_self = CsrAccessPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_valid = early0_EnvPlugin_logic_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_uopId = early0_EnvPlugin_logic_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_4_payload_self = early0_EnvPlugin_logic_flushPort_payload_self;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_valid = DecoderPlugin_logic_laneLogic_0_flushPort_valid;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_uopId = DecoderPlugin_logic_laneLogic_0_flushPort_payload_uopId;
  assign WhiteboxerPlugin_logic_reschedules_flushes_5_payload_self = DecoderPlugin_logic_laneLogic_0_flushPort_payload_self;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_valid = early0_BranchPlugin_logic_jumpLogic_learn_valid;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice = early0_BranchPlugin_logic_jumpLogic_learn_payload_pcOnLastSlice;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget = early0_BranchPlugin_logic_jumpLogic_learn_payload_pcTarget;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken = early0_BranchPlugin_logic_jumpLogic_learn_payload_taken;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch = early0_BranchPlugin_logic_jumpLogic_learn_payload_isBranch;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush = early0_BranchPlugin_logic_jumpLogic_learn_payload_isPush;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop = early0_BranchPlugin_logic_jumpLogic_learn_payload_isPop;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong = early0_BranchPlugin_logic_jumpLogic_learn_payload_wasWrong;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget = early0_BranchPlugin_logic_jumpLogic_learn_payload_badPredictedTarget;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history = early0_BranchPlugin_logic_jumpLogic_learn_payload_history;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId = early0_BranchPlugin_logic_jumpLogic_learn_payload_uopId;
  assign early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = early0_BranchPlugin_logic_jumpLogic_learn_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign WhiteboxerPlugin_logic_prediction_learns_0_valid = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_valid;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_pcOnLastSlice = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcOnLastSlice;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_pcTarget = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_pcTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_taken = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_taken;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isBranch = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isBranch;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isPush = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPush;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_isPop = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_isPop;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_wasWrong = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_wasWrong;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_badPredictedTarget = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_badPredictedTarget;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_history = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_history;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_uopId = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_uopId;
  assign WhiteboxerPlugin_logic_prediction_learns_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = early0_BranchPlugin_logic_jumpLogic_learn_asFlow_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign WhiteboxerPlugin_logic_loadExecute_fire = (((((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && execute_ctrl4_down_AguPlugin_LOAD_lane0) && (! execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0)) && (! execute_ctrl4_down_TRAP_lane0)) && (! execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0));
  assign WhiteboxerPlugin_logic_loadExecute_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_size = execute_ctrl4_down_AguPlugin_SIZE_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_address = execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign WhiteboxerPlugin_logic_loadExecute_data = lane0_IntFormatPlugin_logic_stages_1_wb_payload;
  assign WhiteboxerPlugin_logic_storeCommit_fire = LsuPlugin_logic_onWb_storeFire;
  assign WhiteboxerPlugin_logic_storeCommit_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_size = execute_ctrl4_down_AguPlugin_SIZE_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_address = execute_ctrl4_down_MMU_TRANSLATED_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_data = execute_ctrl4_down_LsuL1_WRITE_DATA_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_storeId = execute_ctrl4_down_Decode_STORE_ID_lane0;
  assign WhiteboxerPlugin_logic_storeCommit_amo = 1'b0;
  assign WhiteboxerPlugin_logic_storeConditional_fire = (((((execute_ctrl4_down_LANE_SEL_lane0 && execute_ctrl4_down_isReady) && (! execute_lane0_ctrls_4_downIsCancel)) && execute_ctrl4_down_AguPlugin_SEL_lane0) && (execute_ctrl4_down_AguPlugin_ATOMIC_lane0 && (! execute_ctrl4_down_AguPlugin_LOAD_lane0))) && (! execute_ctrl4_down_TRAP_lane0));
  assign WhiteboxerPlugin_logic_storeConditional_uopId = execute_ctrl4_down_Decode_UOP_ID_lane0;
  assign WhiteboxerPlugin_logic_storeConditional_miss = execute_ctrl4_down_LsuPlugin_logic_onCtrl_SC_MISS_lane0;
  assign WhiteboxerPlugin_logic_storeBroadcast_fire = LsuPlugin_logic_onWb_storeBroadcast;
  assign WhiteboxerPlugin_logic_storeBroadcast_storeId = execute_ctrl4_down_Decode_STORE_ID_lane0;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_valid = (|lane0_integer_WriteBackPlugin_logic_write_port_valid);
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_address = lane0_integer_WriteBackPlugin_logic_write_port_address;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_data = lane0_integer_WriteBackPlugin_logic_write_port_data;
  assign integer_RegFilePlugin_logic_writeMerges_0_bus_uopId = lane0_integer_WriteBackPlugin_logic_write_port_uopId;
  assign execute_lane0_bypasser_integer_RS1_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_0_data;
  assign execute_lane0_bypasser_integer_RS2_port_data = integer_RegFilePlugin_logic_regfile_fpga_io_reads_1_data;
  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
    if(when_RegFilePlugin_l130) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_valid = 1'b1;
    end
  end

  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
    if(when_RegFilePlugin_l130) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_address = integer_RegFilePlugin_logic_initalizer_counter[4:0];
    end
  end

  always @(*) begin
    integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
    if(when_RegFilePlugin_l130) begin
      integer_RegFilePlugin_logic_regfile_fpga_io_writes_0_data = 32'h0;
    end
  end

  assign integer_RegFilePlugin_logic_initalizer_done = integer_RegFilePlugin_logic_initalizer_counter[5];
  assign when_RegFilePlugin_l130 = (! integer_RegFilePlugin_logic_initalizer_done);
  assign integer_write_0_valid = integer_RegFilePlugin_logic_writeMerges_0_bus_valid;
  assign integer_write_0_address = integer_RegFilePlugin_logic_writeMerges_0_bus_address;
  assign integer_write_0_data = integer_RegFilePlugin_logic_writeMerges_0_bus_data;
  assign integer_write_0_uopId = integer_RegFilePlugin_logic_writeMerges_0_bus_uopId;
  assign execute_freeze_valid = (|{CsrAccessPlugin_logic_fsm_inject_freeze,{LsuPlugin_logic_onCtrl_rva_freezeIt,{LsuPlugin_logic_onCtrl_io_freezeIt,{CfuPlugin_logic_onJoin_freezeIt,{early0_DivPlugin_logic_processing_freeze,CfuPlugin_logic_onFork_freezeIt}}}}});
  assign execute_ctrl5_down_ready = (! execute_freeze_valid);
  assign TrapPlugin_logic_initHold = (|{(! CsrRamPlugin_logic_flush_done),{((! LsuL1Plugin_logic_initializer_done) || 1'b0),{(! integer_RegFilePlugin_logic_initalizer_done),{(FetchL1Plugin_logic_invalidate_firstEver || 1'b0),{1'b0,1'b0}}}}});
  assign WhiteboxerPlugin_logic_wfi = TrapPlugin_logic_harts_0_trap_fsm_wfi;
  assign WhiteboxerPlugin_logic_perf_executeFreezed = execute_freeze_valid;
  assign WhiteboxerPlugin_logic_perf_dispatchHazards = (|(DispatchPlugin_logic_candidates_0_ctx_valid && (! DispatchPlugin_logic_candidates_0_fire)));
  assign WhiteboxerPlugin_logic_perf_candidatesCount = _zz_WhiteboxerPlugin_logic_perf_candidatesCount;
  assign WhiteboxerPlugin_logic_perf_dispatchFeedCount = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCount;
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter = 1'b0;
    if(WhiteboxerPlugin_logic_perf_executeFreezed) begin
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = (_zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 + _zz__zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_executeFreezedCounter = _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2;
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = 1'b0;
    if(WhiteboxerPlugin_logic_perf_dispatchHazards) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchHazardsCounter = _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2;
  assign when_Utils_l586 = (WhiteboxerPlugin_logic_perf_candidatesCount == 1'b0);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = 1'b0;
    if(when_Utils_l586) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_0 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2;
  assign when_Utils_l586_1 = (WhiteboxerPlugin_logic_perf_candidatesCount == 1'b1);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = 1'b0;
    if(when_Utils_l586_1) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = (_zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 + _zz__zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_candidatesCountCounters_1 = _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2;
  assign when_Utils_l586_2 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 1'b0);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = 1'b0;
    if(when_Utils_l586_2) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2;
  assign when_Utils_l586_3 = (WhiteboxerPlugin_logic_perf_dispatchFeedCount == 1'b1);
  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = 1'b0;
    if(when_Utils_l586_3) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = (_zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 + _zz__zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1);
    if(1'b0) begin
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1 = 60'h0;
    end
  end

  assign WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1 = _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2;
  assign WhiteboxerPlugin_logic_trap_ports_0_valid = TrapPlugin_logic_harts_0_trap_whitebox_trap;
  assign WhiteboxerPlugin_logic_trap_ports_0_interrupt = TrapPlugin_logic_harts_0_trap_whitebox_interrupt;
  assign WhiteboxerPlugin_logic_trap_ports_0_cause = TrapPlugin_logic_harts_0_trap_whitebox_code;
  assign fetch_logic_ctrls_2_up_forgetOne = (|fetch_logic_ctrls_2_forgetsSingleRequest_FetchPipelinePlugin_l50);
  assign fetch_logic_ctrls_2_up_cancel = (|fetch_logic_flushes_1_doIt);
  assign fetch_logic_ctrls_1_up_forgetOne = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48);
  assign fetch_logic_ctrls_1_up_cancel = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48);
  assign fetch_logic_ctrls_0_down_ready = fetch_logic_ctrls_1_up_ready;
  assign fetch_logic_ctrls_1_down_ready = fetch_logic_ctrls_2_up_ready;
  always @(*) begin
    fetch_logic_ctrls_0_down_valid = fetch_logic_ctrls_0_up_valid;
    if(when_CtrlLink_l150) begin
      fetch_logic_ctrls_0_down_valid = 1'b0;
    end
  end

  always @(*) begin
    fetch_logic_ctrls_0_up_ready = fetch_logic_ctrls_0_down_isReady;
    if(when_CtrlLink_l150) begin
      fetch_logic_ctrls_0_up_ready = 1'b0;
    end
  end

  assign when_CtrlLink_l150 = (|{fetch_logic_ctrls_0_haltRequest_PcPlugin_l133,{fetch_logic_ctrls_0_haltRequest_BtbPlugin_l200,{fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l297,fetch_logic_ctrls_0_haltRequest_FetchL1Plugin_l217}}});
  assign fetch_logic_ctrls_0_down_Fetch_WORD_PC = fetch_logic_ctrls_0_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_0_down_Fetch_PC_FAULT = fetch_logic_ctrls_0_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_0_down_Fetch_ID = fetch_logic_ctrls_0_up_Fetch_ID;
  always @(*) begin
    fetch_logic_ctrls_1_down_valid = fetch_logic_ctrls_1_up_valid;
    if(when_CtrlLink_l157) begin
      fetch_logic_ctrls_1_down_valid = 1'b0;
    end
  end

  assign fetch_logic_ctrls_1_up_ready = fetch_logic_ctrls_1_down_isReady;
  assign when_CtrlLink_l157 = (|fetch_logic_ctrls_1_throwWhen_FetchPipelinePlugin_l48);
  assign fetch_logic_ctrls_1_down_Fetch_WORD_PC = fetch_logic_ctrls_1_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_1_down_Fetch_PC_FAULT = fetch_logic_ctrls_1_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_1_down_Fetch_ID = fetch_logic_ctrls_1_up_Fetch_ID;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_1 = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_1;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
  assign fetch_logic_ctrls_1_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS = fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_HASH = fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH;
  assign fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY = fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_valid = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_address = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address;
  assign fetch_logic_ctrls_1_down_GSharePlugin_logic_BYPASS_payload_data_0 = fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0;
  assign fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS = fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS;
  assign fetch_logic_ctrls_2_down_valid = fetch_logic_ctrls_2_up_valid;
  assign fetch_logic_ctrls_2_up_ready = fetch_logic_ctrls_2_down_isReady;
  assign fetch_logic_ctrls_2_down_Fetch_WORD_PC = fetch_logic_ctrls_2_up_Fetch_WORD_PC;
  assign fetch_logic_ctrls_2_down_Fetch_PC_FAULT = fetch_logic_ctrls_2_up_Fetch_PC_FAULT;
  assign fetch_logic_ctrls_2_down_Fetch_ID = fetch_logic_ctrls_2_up_Fetch_ID;
  assign fetch_logic_ctrls_2_down_Prediction_BRANCH_HISTORY = fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_0_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_1_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_2_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_2_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_2_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_2_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_2_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_2_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_3_loaded = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_3_loaded;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_3_error = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_3_error;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_TAGS_3_address = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_3_address;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_PLRU_BYPASSED_1 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_1;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_1 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_2 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_2;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_BANKS_MUXES_3 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_3;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_HAZARD = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_0 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_1 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_2 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_2;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HITS_3 = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_3;
  assign fetch_logic_ctrls_2_down_MMU_BYPASS_TRANSLATION = fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION;
  assign fetch_logic_ctrls_2_down_FetchL1Plugin_logic_WAYS_HIT = fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT;
  assign fetch_logic_ctrls_2_down_GSharePlugin_GSHARE_COUNTER_0 = fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMPED = fetch_logic_ctrls_2_up_Prediction_WORD_JUMPED;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_JUMP_PC = fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_PC;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_BRANCH = fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_BRANCH;
  assign fetch_logic_ctrls_2_down_Prediction_WORD_SLICES_TAKEN = fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_TAKEN;
  assign fetch_logic_ctrls_2_down_MMU_HAZARD = fetch_logic_ctrls_2_up_MMU_HAZARD;
  assign fetch_logic_ctrls_2_down_MMU_REFILL = fetch_logic_ctrls_2_up_MMU_REFILL;
  assign fetch_logic_ctrls_2_down_MMU_TRANSLATED = fetch_logic_ctrls_2_up_MMU_TRANSLATED;
  assign fetch_logic_ctrls_2_down_MMU_ALLOW_EXECUTE = fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE;
  assign fetch_logic_ctrls_2_down_MMU_PAGE_FAULT = fetch_logic_ctrls_2_up_MMU_PAGE_FAULT;
  assign fetch_logic_ctrls_2_down_MMU_ACCESS_FAULT = fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT;
  always @(*) begin
    decode_ctrls_0_down_ready = decode_ctrls_1_up_ready;
    if(when_StageLink_l67) begin
      decode_ctrls_0_down_ready = 1'b1;
    end
  end

  assign when_StageLink_l67 = (! decode_ctrls_1_up_isValid);
  assign when_DecodePipelinePlugin_l70 = ((! decode_ctrls_1_up_isReady) && decode_ctrls_1_lane0_upIsCancel);
  assign decode_ctrls_0_down_valid = decode_ctrls_0_up_valid;
  assign decode_ctrls_0_up_ready = decode_ctrls_0_down_isReady;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_0 = decode_ctrls_0_up_Decode_INSTRUCTION_0;
  assign decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0 = decode_ctrls_0_up_Decode_DECOMPRESSION_FAULT_0;
  assign decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0 = decode_ctrls_0_up_Decode_INSTRUCTION_RAW_0;
  assign decode_ctrls_0_down_PC_0 = decode_ctrls_0_up_PC_0;
  assign decode_ctrls_0_down_Decode_DOP_ID_0 = decode_ctrls_0_up_Decode_DOP_ID_0;
  assign decode_ctrls_0_down_Fetch_ID_0 = decode_ctrls_0_up_Fetch_ID_0;
  assign decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0 = decode_ctrls_0_up_GSharePlugin_GSHARE_COUNTER_0_0;
  assign decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0 = decode_ctrls_0_up_Prediction_BRANCH_HISTORY_0;
  assign decode_ctrls_0_down_TRAP_0 = decode_ctrls_0_up_TRAP_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0 = decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0 = decode_ctrls_0_up_Prediction_ALIGNED_JUMPED_PC_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0 = decode_ctrls_0_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0 = decode_ctrls_0_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign decode_ctrls_0_down_Prediction_ALIGN_REDO_0 = decode_ctrls_0_up_Prediction_ALIGN_REDO_0;
  assign decode_ctrls_1_down_valid = decode_ctrls_1_up_valid;
  assign decode_ctrls_1_up_ready = decode_ctrls_1_down_isReady;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_0 = decode_ctrls_1_up_Decode_INSTRUCTION_0;
  assign decode_ctrls_1_down_Decode_DECOMPRESSION_FAULT_0 = decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0;
  assign decode_ctrls_1_down_Decode_INSTRUCTION_RAW_0 = decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0;
  assign decode_ctrls_1_down_PC_0 = decode_ctrls_1_up_PC_0;
  assign decode_ctrls_1_down_Decode_DOP_ID_0 = decode_ctrls_1_up_Decode_DOP_ID_0;
  assign decode_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0_0 = decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0;
  assign decode_ctrls_1_down_Prediction_BRANCH_HISTORY_0 = decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_0 = decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_JUMPED_PC_0 = decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_SLICES_BRANCH_0 = decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0;
  assign decode_ctrls_1_down_Prediction_ALIGNED_SLICES_TAKEN_0 = decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0;
  assign decode_ctrls_1_down_Prediction_ALIGN_REDO_0 = decode_ctrls_1_up_Prediction_ALIGN_REDO_0;
  assign execute_ctrl0_down_ready = execute_ctrl1_up_ready;
  assign execute_ctrl1_down_ready = execute_ctrl2_up_ready;
  assign execute_ctrl2_down_ready = execute_ctrl3_up_ready;
  assign execute_ctrl3_down_ready = execute_ctrl4_up_ready;
  assign execute_ctrl4_down_ready = execute_ctrl5_up_ready;
  assign execute_ctrl0_up_ready = execute_ctrl0_down_isReady;
  assign execute_ctrl0_down_Decode_UOP_lane0 = execute_ctrl0_up_Decode_UOP_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl0_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl0_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl0_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl0_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl0_down_PC_lane0 = execute_ctrl0_up_PC_lane0;
  assign execute_ctrl0_down_TRAP_lane0 = execute_ctrl0_up_TRAP_lane0;
  assign execute_ctrl0_down_Decode_UOP_ID_lane0 = execute_ctrl0_up_Decode_UOP_ID_lane0;
  assign execute_ctrl0_down_RS1_PHYS_lane0 = execute_ctrl0_up_RS1_PHYS_lane0;
  assign execute_ctrl0_down_RS2_PHYS_lane0 = execute_ctrl0_up_RS2_PHYS_lane0;
  assign execute_ctrl0_down_RD_PHYS_lane0 = execute_ctrl0_up_RD_PHYS_lane0;
  assign execute_ctrl0_down_COMPLETED_lane0 = execute_ctrl0_up_COMPLETED_lane0;
  assign execute_ctrl1_up_ready = execute_ctrl1_down_isReady;
  assign execute_ctrl1_down_Decode_UOP_lane0 = execute_ctrl1_up_Decode_UOP_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl1_down_PC_lane0 = execute_ctrl1_up_PC_lane0;
  assign execute_ctrl1_down_TRAP_lane0 = execute_ctrl1_up_TRAP_lane0;
  assign execute_ctrl1_down_Decode_UOP_ID_lane0 = execute_ctrl1_up_Decode_UOP_ID_lane0;
  assign execute_ctrl1_down_RS1_PHYS_lane0 = execute_ctrl1_up_RS1_PHYS_lane0;
  assign execute_ctrl1_down_RS2_PHYS_lane0 = execute_ctrl1_up_RS2_PHYS_lane0;
  assign execute_ctrl1_down_RD_PHYS_lane0 = execute_ctrl1_up_RD_PHYS_lane0;
  assign execute_ctrl1_down_COMPLETED_lane0 = execute_ctrl1_up_COMPLETED_lane0;
  assign execute_ctrl1_down_AguPlugin_SIZE_lane0 = execute_ctrl1_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl2_up_ready = execute_ctrl2_down_isReady;
  assign execute_ctrl2_down_Decode_UOP_lane0 = execute_ctrl2_up_Decode_UOP_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl2_down_Prediction_ALIGNED_JUMPED_PC_lane0 = execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0;
  assign execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl2_down_PC_lane0 = execute_ctrl2_up_PC_lane0;
  assign execute_ctrl2_down_Decode_UOP_ID_lane0 = execute_ctrl2_up_Decode_UOP_ID_lane0;
  assign execute_ctrl2_down_RD_PHYS_lane0 = execute_ctrl2_up_RD_PHYS_lane0;
  assign execute_ctrl2_down_AguPlugin_SIZE_lane0 = execute_ctrl2_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl2_down_early0_SrcPlugin_SRC1_lane0 = execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0;
  assign execute_ctrl2_down_early0_SrcPlugin_SRC2_lane0 = execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0;
  assign execute_ctrl2_down_integer_RS2_lane0 = execute_ctrl2_up_integer_RS2_lane0;
  assign execute_ctrl2_down_MAY_FLUSH_PRECISE_3_lane0 = execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_SEL_lane0 = execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_BarrelShifterPlugin_SEL_lane0 = execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_BranchPlugin_SEL_lane0 = execute_ctrl2_up_early0_BranchPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_MulPlugin_SEL_lane0 = execute_ctrl2_up_early0_MulPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_DivPlugin_SEL_lane0 = execute_ctrl2_up_early0_DivPlugin_SEL_lane0;
  assign execute_ctrl2_down_early0_EnvPlugin_SEL_lane0 = execute_ctrl2_up_early0_EnvPlugin_SEL_lane0;
  assign execute_ctrl2_down_CfuPlugin_logic_CFU_ENABLE_lane0 = execute_ctrl2_up_CfuPlugin_logic_CFU_ENABLE_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 = execute_ctrl2_up_CsrAccessPlugin_SEL_lane0;
  assign execute_ctrl2_down_AguPlugin_SEL_lane0 = execute_ctrl2_up_AguPlugin_SEL_lane0;
  assign execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0 = execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0;
  assign execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0 = execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_2_lane0 = execute_ctrl2_up_COMPLETION_AT_2_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_3_lane0 = execute_ctrl2_up_COMPLETION_AT_3_lane0;
  assign execute_ctrl2_down_COMPLETION_AT_4_lane0 = execute_ctrl2_up_COMPLETION_AT_4_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl2_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl2_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0 = execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_SLTX_lane0 = execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0;
  assign execute_ctrl2_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 = execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
  assign execute_ctrl2_down_SrcStageables_REVERT_lane0 = execute_ctrl2_up_SrcStageables_REVERT_lane0;
  assign execute_ctrl2_down_SrcStageables_ZERO_lane0 = execute_ctrl2_up_SrcStageables_ZERO_lane0;
  assign execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign execute_ctrl2_down_BYPASSED_AT_3_lane0 = execute_ctrl2_up_BYPASSED_AT_3_lane0;
  assign execute_ctrl2_down_SrcStageables_UNSIGNED_lane0 = execute_ctrl2_up_SrcStageables_UNSIGNED_lane0;
  assign execute_ctrl2_down_BarrelShifterPlugin_LEFT_lane0 = execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0;
  assign execute_ctrl2_down_BarrelShifterPlugin_SIGNED_lane0 = execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0;
  assign execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0 = execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0;
  assign execute_ctrl2_down_CfuPlugin_logic_CFU_ENCODING_lane0 = execute_ctrl2_up_CfuPlugin_logic_CFU_ENCODING_lane0;
  assign execute_ctrl2_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0 = execute_ctrl2_up_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0;
  assign execute_ctrl2_down_MulPlugin_HIGH_lane0 = execute_ctrl2_up_MulPlugin_HIGH_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS1_SIGNED_lane0 = execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0;
  assign execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0 = execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0;
  assign execute_ctrl2_down_DivPlugin_REM_lane0 = execute_ctrl2_up_DivPlugin_REM_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_CSR_IMM_lane0 = execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_CSR_MASK_lane0 = execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0;
  assign execute_ctrl2_down_CsrAccessPlugin_CSR_CLEAR_lane0 = execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0;
  assign execute_ctrl2_down_AguPlugin_LOAD_lane0 = execute_ctrl2_up_AguPlugin_LOAD_lane0;
  assign execute_ctrl2_down_AguPlugin_STORE_lane0 = execute_ctrl2_up_AguPlugin_STORE_lane0;
  assign execute_ctrl2_down_AguPlugin_ATOMIC_lane0 = execute_ctrl2_up_AguPlugin_ATOMIC_lane0;
  assign execute_ctrl2_down_AguPlugin_FLOAT_lane0 = execute_ctrl2_up_AguPlugin_FLOAT_lane0;
  assign execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign execute_ctrl2_down_early0_EnvPlugin_OP_lane0 = execute_ctrl2_up_early0_EnvPlugin_OP_lane0;
  assign execute_ctrl3_up_ready = execute_ctrl3_down_isReady;
  assign execute_ctrl3_down_Decode_UOP_lane0 = execute_ctrl3_up_Decode_UOP_lane0;
  assign execute_ctrl3_down_Prediction_ALIGNED_JUMPED_lane0 = execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane0;
  assign execute_ctrl3_down_GSharePlugin_GSHARE_COUNTER_lane0_0 = execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_0;
  assign execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl3_down_PC_lane0 = execute_ctrl3_up_PC_lane0;
  assign execute_ctrl3_down_Decode_UOP_ID_lane0 = execute_ctrl3_up_Decode_UOP_ID_lane0;
  assign execute_ctrl3_down_RD_PHYS_lane0 = execute_ctrl3_up_RD_PHYS_lane0;
  assign execute_ctrl3_down_AguPlugin_SIZE_lane0 = execute_ctrl3_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl3_down_integer_RS2_lane0 = execute_ctrl3_up_integer_RS2_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_SEL_lane0 = execute_ctrl3_up_early0_BranchPlugin_SEL_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_SEL_lane0 = execute_ctrl3_up_early0_MulPlugin_SEL_lane0;
  assign execute_ctrl3_down_early0_DivPlugin_SEL_lane0 = execute_ctrl3_up_early0_DivPlugin_SEL_lane0;
  assign execute_ctrl3_down_CfuPlugin_logic_CFU_ENABLE_lane0 = execute_ctrl3_up_CfuPlugin_logic_CFU_ENABLE_lane0;
  assign execute_ctrl3_down_CsrAccessPlugin_SEL_lane0 = execute_ctrl3_up_CsrAccessPlugin_SEL_lane0;
  assign execute_ctrl3_down_AguPlugin_SEL_lane0 = execute_ctrl3_up_AguPlugin_SEL_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0 = execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0;
  assign execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0 = execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_3_lane0 = execute_ctrl3_up_COMPLETION_AT_3_lane0;
  assign execute_ctrl3_down_COMPLETION_AT_4_lane0 = execute_ctrl3_up_COMPLETION_AT_4_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
  assign execute_ctrl3_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl3_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign execute_ctrl3_down_BranchPlugin_BRANCH_CTRL_lane0 = execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0;
  assign execute_ctrl3_down_MulPlugin_HIGH_lane0 = execute_ctrl3_up_MulPlugin_HIGH_lane0;
  assign execute_ctrl3_down_AguPlugin_LOAD_lane0 = execute_ctrl3_up_AguPlugin_LOAD_lane0;
  assign execute_ctrl3_down_AguPlugin_STORE_lane0 = execute_ctrl3_up_AguPlugin_STORE_lane0;
  assign execute_ctrl3_down_AguPlugin_ATOMIC_lane0 = execute_ctrl3_up_AguPlugin_ATOMIC_lane0;
  assign execute_ctrl3_down_AguPlugin_FLOAT_lane0 = execute_ctrl3_up_AguPlugin_FLOAT_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign execute_ctrl3_down_early0_SrcPlugin_ADD_SUB_lane0 = execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0;
  assign execute_ctrl3_down_early0_SrcPlugin_LESS_lane0 = execute_ctrl3_up_early0_SrcPlugin_LESS_lane0;
  assign execute_ctrl3_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0 = execute_ctrl3_up_CfuPlugin_logic_CFU_IN_FLIGHT_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  assign execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  assign execute_ctrl3_down_DivPlugin_DIV_RESULT_lane0 = execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 = execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 = execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 = execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_logic_alu_EQ_lane0 = execute_ctrl3_up_early0_BranchPlugin_logic_alu_EQ_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 = execute_ctrl3_up_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
  assign execute_ctrl3_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 = execute_ctrl3_up_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
  assign execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0 = execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_1 = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_1;
  assign execute_ctrl3_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty = execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  assign execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0 = execute_ctrl3_up_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  assign execute_ctrl3_down_LsuL1_MASK_lane0 = execute_ctrl3_up_LsuL1_MASK_lane0;
  assign execute_ctrl3_down_LsuL1_SIZE_lane0 = execute_ctrl3_up_LsuL1_SIZE_lane0;
  assign execute_ctrl3_down_LsuL1_LOAD_lane0 = execute_ctrl3_up_LsuL1_LOAD_lane0;
  assign execute_ctrl3_down_LsuL1_ATOMIC_lane0 = execute_ctrl3_up_LsuL1_ATOMIC_lane0;
  assign execute_ctrl3_down_LsuL1_STORE_lane0 = execute_ctrl3_up_LsuL1_STORE_lane0;
  assign execute_ctrl3_down_LsuL1_CLEAN_lane0 = execute_ctrl3_up_LsuL1_CLEAN_lane0;
  assign execute_ctrl3_down_LsuL1_INVALID_lane0 = execute_ctrl3_up_LsuL1_INVALID_lane0;
  assign execute_ctrl3_down_LsuL1_PREFETCH_lane0 = execute_ctrl3_up_LsuL1_PREFETCH_lane0;
  assign execute_ctrl3_down_LsuL1_FLUSH_lane0 = execute_ctrl3_up_LsuL1_FLUSH_lane0;
  assign execute_ctrl3_down_Decode_STORE_ID_lane0 = execute_ctrl3_up_Decode_STORE_ID_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0;
  assign execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_valid = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_valid;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_virtualAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_virtualAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_physicalAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_physicalAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowRead = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowRead;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowWrite = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowWrite;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowExecute = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowExecute;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_0_allowUser = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowUser;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_valid = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_valid;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_virtualAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_virtualAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_physicalAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_physicalAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowRead = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowRead;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowWrite = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowWrite;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowExecute = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowExecute;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_1_allowUser = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowUser;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_valid = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_valid;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_virtualAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_virtualAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_physicalAddress = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_physicalAddress;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowRead = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowRead;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowWrite = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowWrite;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowExecute = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowExecute;
  assign execute_ctrl3_down_MMU_L0_ENTRIES_lane0_2_allowUser = execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowUser;
  assign execute_ctrl3_down_MMU_L0_HITS_PRE_VALID_lane0 = execute_ctrl3_up_MMU_L0_HITS_PRE_VALID_lane0;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_valid = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_valid;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_virtualAddress = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_virtualAddress;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_physicalAddress = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_physicalAddress;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowRead = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowRead;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowWrite = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowWrite;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowExecute = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowExecute;
  assign execute_ctrl3_down_MMU_L1_ENTRIES_lane0_0_allowUser = execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowUser;
  assign execute_ctrl3_down_MMU_L1_HITS_PRE_VALID_lane0 = execute_ctrl3_up_MMU_L1_HITS_PRE_VALID_lane0;
  assign execute_ctrl4_up_ready = execute_ctrl4_down_isReady;
  assign execute_ctrl4_down_Decode_UOP_lane0 = execute_ctrl4_up_Decode_UOP_lane0;
  assign execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0 = execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0;
  assign execute_ctrl4_down_PC_lane0 = execute_ctrl4_up_PC_lane0;
  assign execute_ctrl4_down_Decode_UOP_ID_lane0 = execute_ctrl4_up_Decode_UOP_ID_lane0;
  assign execute_ctrl4_down_RD_PHYS_lane0 = execute_ctrl4_up_RD_PHYS_lane0;
  assign execute_ctrl4_down_AguPlugin_SIZE_lane0 = execute_ctrl4_up_AguPlugin_SIZE_lane0;
  assign execute_ctrl4_down_integer_RS2_lane0 = execute_ctrl4_up_integer_RS2_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_SEL_lane0 = execute_ctrl4_up_early0_MulPlugin_SEL_lane0;
  assign execute_ctrl4_down_CfuPlugin_logic_CFU_ENABLE_lane0 = execute_ctrl4_up_CfuPlugin_logic_CFU_ENABLE_lane0;
  assign execute_ctrl4_down_AguPlugin_SEL_lane0 = execute_ctrl4_up_AguPlugin_SEL_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FENCE_lane0 = execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0;
  assign execute_ctrl4_down_lane0_integer_WriteBackPlugin_SEL_lane0 = execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0;
  assign execute_ctrl4_down_COMPLETION_AT_4_lane0 = execute_ctrl4_up_COMPLETION_AT_4_lane0;
  assign execute_ctrl4_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0 = execute_ctrl4_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
  assign execute_ctrl4_down_lane0_IntFormatPlugin_logic_SIGNED_lane0 = execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0;
  assign execute_ctrl4_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 = execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
  assign execute_ctrl4_down_MulPlugin_HIGH_lane0 = execute_ctrl4_up_MulPlugin_HIGH_lane0;
  assign execute_ctrl4_down_AguPlugin_LOAD_lane0 = execute_ctrl4_up_AguPlugin_LOAD_lane0;
  assign execute_ctrl4_down_AguPlugin_STORE_lane0 = execute_ctrl4_up_AguPlugin_STORE_lane0;
  assign execute_ctrl4_down_AguPlugin_ATOMIC_lane0 = execute_ctrl4_up_AguPlugin_ATOMIC_lane0;
  assign execute_ctrl4_down_AguPlugin_FLOAT_lane0 = execute_ctrl4_up_AguPlugin_FLOAT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_LSU_PREFETCH_lane0 = execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0;
  assign execute_ctrl4_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0 = execute_ctrl4_up_CfuPlugin_logic_CFU_IN_FLIGHT_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_0_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_0_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_1_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_1_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_2_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_2_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_mul_VALUES_3_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_3_lane0;
  assign execute_ctrl4_down_LsuL1_MIXED_ADDRESS_lane0 = execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FROM_ACCESS_lane0 = execute_ctrl4_up_LsuPlugin_logic_FROM_ACCESS_lane0;
  assign execute_ctrl4_down_LsuL1_MASK_lane0 = execute_ctrl4_up_LsuL1_MASK_lane0;
  assign execute_ctrl4_down_LsuL1_SIZE_lane0 = execute_ctrl4_up_LsuL1_SIZE_lane0;
  assign execute_ctrl4_down_LsuL1_LOAD_lane0 = execute_ctrl4_up_LsuL1_LOAD_lane0;
  assign execute_ctrl4_down_LsuL1_ATOMIC_lane0 = execute_ctrl4_up_LsuL1_ATOMIC_lane0;
  assign execute_ctrl4_down_LsuL1_STORE_lane0 = execute_ctrl4_up_LsuL1_STORE_lane0;
  assign execute_ctrl4_down_LsuL1_CLEAN_lane0 = execute_ctrl4_up_LsuL1_CLEAN_lane0;
  assign execute_ctrl4_down_LsuL1_INVALID_lane0 = execute_ctrl4_up_LsuL1_INVALID_lane0;
  assign execute_ctrl4_down_LsuL1_PREFETCH_lane0 = execute_ctrl4_up_LsuL1_PREFETCH_lane0;
  assign execute_ctrl4_down_LsuL1_FLUSH_lane0 = execute_ctrl4_up_LsuL1_FLUSH_lane0;
  assign execute_ctrl4_down_Decode_STORE_ID_lane0 = execute_ctrl4_up_Decode_STORE_ID_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FROM_LSU_lane0 = execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_FROM_PREFETCH_lane0 = execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_0 = execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_plru_1 = execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_1;
  assign execute_ctrl4_down_LsuL1Plugin_logic_SHARED_lane0_dirty = execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty;
  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_0_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0;
  assign execute_ctrl4_down_early0_MulPlugin_logic_steps_0_adders_1_lane0 = execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 = execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 = execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2 = execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_2;
  assign execute_ctrl4_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3 = execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_3;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
  assign execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0 = execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault;
  assign execute_ctrl4_down_LsuL1Plugin_logic_WAYS_HITS_lane0 = execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onTrigger_HIT_lane0 = execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0;
  assign execute_ctrl4_down_MMU_TRANSLATED_lane0 = execute_ctrl4_up_MMU_TRANSLATED_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 = execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0 = execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault = execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io = execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault = execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io = execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_IO_lane0 = execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 = execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 = execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
  assign execute_ctrl4_down_LsuPlugin_logic_MMU_FAILURE_lane0 = execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0;
  assign execute_ctrl4_down_MMU_ACCESS_FAULT_lane0 = execute_ctrl4_up_MMU_ACCESS_FAULT_lane0;
  assign execute_ctrl4_down_MMU_REFILL_lane0 = execute_ctrl4_up_MMU_REFILL_lane0;
  assign execute_ctrl4_down_MMU_HAZARD_lane0 = execute_ctrl4_up_MMU_HAZARD_lane0;
  assign execute_ctrl4_down_MMU_BYPASS_TRANSLATION_lane0 = execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0;
  assign execute_ctrl5_up_ready = execute_ctrl5_down_isReady;
  assign execute_ctrl5_down_LANE_SEL_lane0 = execute_ctrl5_up_LANE_SEL_lane0;
  assign execute_ctrl5_down_RD_PHYS_lane0 = execute_ctrl5_up_RD_PHYS_lane0;
  assign execute_ctrl5_down_COMMIT_lane0 = execute_ctrl5_up_COMMIT_lane0;
  assign execute_ctrl5_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0 = execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
  assign fetch_logic_ctrls_0_down_isFiring = (fetch_logic_ctrls_0_down_isValid && fetch_logic_ctrls_0_down_isReady);
  assign fetch_logic_ctrls_0_down_isValid = fetch_logic_ctrls_0_down_valid;
  assign fetch_logic_ctrls_0_down_isReady = fetch_logic_ctrls_0_down_ready;
  assign fetch_logic_ctrls_1_up_isValid = fetch_logic_ctrls_1_up_valid;
  assign fetch_logic_ctrls_1_up_isReady = fetch_logic_ctrls_1_up_ready;
  assign fetch_logic_ctrls_1_up_isCancel = fetch_logic_ctrls_1_up_cancel;
  assign fetch_logic_ctrls_1_down_isValid = fetch_logic_ctrls_1_down_valid;
  assign fetch_logic_ctrls_1_down_isReady = fetch_logic_ctrls_1_down_ready;
  assign fetch_logic_ctrls_2_up_isMoving = (fetch_logic_ctrls_2_up_isValid && (fetch_logic_ctrls_2_up_isReady || fetch_logic_ctrls_2_up_isCancel));
  assign fetch_logic_ctrls_2_up_isValid = fetch_logic_ctrls_2_up_valid;
  assign fetch_logic_ctrls_2_up_isReady = fetch_logic_ctrls_2_up_ready;
  assign fetch_logic_ctrls_2_up_isCancel = fetch_logic_ctrls_2_up_cancel;
  assign fetch_logic_ctrls_2_up_isCanceling = (fetch_logic_ctrls_2_up_isValid && fetch_logic_ctrls_2_up_isCancel);
  assign fetch_logic_ctrls_0_up_isFiring = (fetch_logic_ctrls_0_up_isValid && fetch_logic_ctrls_0_up_isReady);
  assign fetch_logic_ctrls_0_up_isValid = fetch_logic_ctrls_0_up_valid;
  assign fetch_logic_ctrls_0_up_isReady = fetch_logic_ctrls_0_up_ready;
  assign fetch_logic_ctrls_2_down_isValid = fetch_logic_ctrls_2_down_valid;
  assign fetch_logic_ctrls_2_down_isReady = fetch_logic_ctrls_2_down_ready;
  assign decode_ctrls_0_down_isValid = decode_ctrls_0_down_valid;
  assign decode_ctrls_0_down_isReady = decode_ctrls_0_down_ready;
  assign decode_ctrls_1_up_isMoving = (decode_ctrls_1_up_isValid && decode_ctrls_1_up_isReady);
  assign decode_ctrls_1_up_isValid = decode_ctrls_1_up_valid;
  assign decode_ctrls_1_up_isReady = decode_ctrls_1_up_ready;
  assign decode_ctrls_1_up_isCanceling = 1'b0;
  assign decode_ctrls_0_up_isFiring = (decode_ctrls_0_up_isValid && decode_ctrls_0_up_isReady);
  assign decode_ctrls_0_up_isMoving = (decode_ctrls_0_up_isValid && decode_ctrls_0_up_isReady);
  assign decode_ctrls_0_up_isValid = decode_ctrls_0_up_valid;
  assign decode_ctrls_0_up_isReady = decode_ctrls_0_up_ready;
  assign decode_ctrls_1_down_isReady = decode_ctrls_1_down_ready;
  assign execute_ctrl0_down_isReady = execute_ctrl0_down_ready;
  assign execute_ctrl1_down_isReady = execute_ctrl1_down_ready;
  assign execute_ctrl2_down_isReady = execute_ctrl2_down_ready;
  assign execute_ctrl3_down_isReady = execute_ctrl3_down_ready;
  assign execute_ctrl4_up_isReady = execute_ctrl4_up_ready;
  assign execute_ctrl4_down_isReady = execute_ctrl4_down_ready;
  assign execute_ctrl5_down_isReady = execute_ctrl5_down_ready;
  always @(*) begin
    LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_stateReg;
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_CMD : begin
        if(when_LsuPlugin_l363) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_COMPLETION;
        end
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
        if(when_LsuPlugin_l371) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_IDLE;
        end
      end
      default : begin
        if(LsuPlugin_logic_flusher_arbiter_io_output_valid) begin
          LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_CMD;
        end
      end
    endcase
    if(LsuPlugin_logic_flusher_wantKill) begin
      LsuPlugin_logic_flusher_stateNext = LsuPlugin_logic_flusher_IDLE;
    end
  end

  assign when_LsuPlugin_l363 = (LsuPlugin_logic_flusher_cmdCounter[6] && (! LsuPlugin_logic_flusher_inflight));
  assign when_LsuPlugin_l371 = (! (|LsuPlugin_logic_flusher_waiter));
  assign LsuPlugin_logic_flusher_onExit_IDLE = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_IDLE) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_IDLE));
  assign LsuPlugin_logic_flusher_onExit_CMD = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_CMD) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_CMD));
  assign LsuPlugin_logic_flusher_onExit_COMPLETION = ((LsuPlugin_logic_flusher_stateNext != LsuPlugin_logic_flusher_COMPLETION) && (LsuPlugin_logic_flusher_stateReg == LsuPlugin_logic_flusher_COMPLETION));
  assign LsuPlugin_logic_flusher_onEntry_IDLE = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_IDLE) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_IDLE));
  assign LsuPlugin_logic_flusher_onEntry_CMD = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_CMD) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_CMD));
  assign LsuPlugin_logic_flusher_onEntry_COMPLETION = ((LsuPlugin_logic_flusher_stateNext == LsuPlugin_logic_flusher_COMPLETION) && (LsuPlugin_logic_flusher_stateReg != LsuPlugin_logic_flusher_COMPLETION));
  always @(*) begin
    TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_stateReg;
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
        if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
        if(when_TrapPlugin_l409) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL;
        end else begin
          case(TrapPlugin_logic_harts_0_trap_pending_state_code)
            4'b0000 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
            end
            4'b0001 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC;
            end
            4'b0010 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH;
            end
            4'b0100 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
            end
            4'b0101 : begin
              TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
            end
            4'b1000 : begin
              if(TrapPlugin_api_harts_0_askWake) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
              end
            end
            4'b0110 : begin
              if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_ready) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
              end
            end
            4'b0111 : begin
              if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_cmd_ready) begin
                TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP;
              end
            end
            default : begin
            end
          endcase
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_write_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        if(TrapPlugin_logic_harts_0_crsPorts_write_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_read_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        if(TrapPlugin_logic_harts_0_crsPorts_read_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
        if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
          if(when_TrapPlugin_l509) begin
            TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL;
          end
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
        if(TrapPlugin_logic_lsuL1Invalidate_0_cmd_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH;
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
        if(TrapPlugin_logic_fetchL1Invalidate_0_cmd_ready) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_JUMP;
        end
      end
      default : begin
        if(when_TrapPlugin_l362) begin
          TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RUNNING;
        end
      end
    endcase
    if(TrapPlugin_logic_harts_0_trap_fsm_wantKill) begin
      TrapPlugin_logic_harts_0_trap_fsm_stateNext = TrapPlugin_logic_harts_0_trap_fsm_RESET;
    end
  end

  assign when_TrapPlugin_l409 = ((TrapPlugin_logic_harts_0_trap_pending_state_exception || TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak) || TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt);
  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address = 4'b1001;
    case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_write_address = 4'b0101;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1 = 4'b1010;
    case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_write_address_1 = 4'b0110;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address = 4'b1011;
    case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_read_address = 4'b0111;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1 = 4'b1001;
    case(TrapPlugin_logic_harts_0_trap_fsm_xretPrivilege)
      2'b01 : begin
        _zz_TrapPlugin_logic_harts_0_crsPorts_read_address_1 = 4'b0101;
      end
      default : begin
      end
    endcase
  end

  assign when_TrapPlugin_l654 = (TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege != 2'b11);
  assign switch_TrapPlugin_l655 = TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0];
  assign when_TrapPlugin_l509 = (TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_pageFault || TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault);
  assign switch_TrapPlugin_l511 = {TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_payload_accessFault,TrapPlugin_logic_harts_0_trap_pending_state_arg[1 : 0]};
  assign when_TrapPlugin_l362 = (&{TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated,TrapPlugin_logic_harts_0_trap_fsm_resetToRunConditions_0});
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_RESET = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_RESET) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RESET));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_RUNNING = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_RUNNING) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_RUNNING));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_PROCESS_1 = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVAL = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_TVEC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_TRAP_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_XRET_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_ATS_RSP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_JUMP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_JUMP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_JUMP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_LSU_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH));
  assign TrapPlugin_logic_harts_0_trap_fsm_onExit_FETCH_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext != TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg == TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_RESET = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_RESET) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_RESET));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_RUNNING = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_RUNNING) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_RUNNING));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_PROCESS_1 = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVAL = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_TVEC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_TRAP_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_EPC = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_XRET_APPLY = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_ATS_RSP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_JUMP = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_JUMP) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_JUMP));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_LSU_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH));
  assign TrapPlugin_logic_harts_0_trap_fsm_onEntry_FETCH_FLUSH = ((TrapPlugin_logic_harts_0_trap_fsm_stateNext == TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH) && (TrapPlugin_logic_harts_0_trap_fsm_stateReg != TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH));
  always @(*) begin
    MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_stateReg;
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
        if(MmuPlugin_logic_refill_arbiter_io_output_valid) begin
          MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_1;
        end
      end
      MmuPlugin_logic_refill_CMD_0 : begin
        if(when_MmuPlugin_l470) begin
          if(MmuPlugin_logic_accessBus_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_RSP_0;
          end
        end
      end
      MmuPlugin_logic_refill_CMD_1 : begin
        if(when_MmuPlugin_l470_1) begin
          if(MmuPlugin_logic_accessBus_cmd_ready) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_RSP_1;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_0 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_0;
          end else begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_IDLE;
          end
        end
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_1;
          end else begin
            if(when_MmuPlugin_l487) begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_IDLE;
            end else begin
              MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_CMD_0;
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(MmuPlugin_logic_refill_wantStart) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_IDLE;
    end
    if(MmuPlugin_logic_refill_wantKill) begin
      MmuPlugin_logic_refill_stateNext = MmuPlugin_logic_refill_BOOT;
    end
  end

  assign when_MmuPlugin_l470 = (1'b1 && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l470_1 = (1'b1 && (MmuPlugin_logic_refill_cacheRefillAny == 1'b0));
  assign when_MmuPlugin_l479 = (! MmuPlugin_logic_refill_load_leaf);
  assign when_MmuPlugin_l455 = (MmuPlugin_logic_refill_fetch_0_pageFault || MmuPlugin_logic_refill_fetch_0_accessFault);
  assign _zz_57 = MmuPlugin_logic_refill_portOhReg[0];
  assign when_MmuPlugin_l455_1 = (MmuPlugin_logic_refill_fetch_0_pageFault || MmuPlugin_logic_refill_fetch_0_accessFault);
  assign when_MmuPlugin_l487 = (MmuPlugin_logic_refill_load_leaf || MmuPlugin_logic_refill_load_exception);
  assign when_MmuPlugin_l455_2 = (MmuPlugin_logic_refill_fetch_1_pageFault || MmuPlugin_logic_refill_fetch_1_accessFault);
  assign when_MmuPlugin_l455_3 = (MmuPlugin_logic_refill_fetch_1_pageFault || MmuPlugin_logic_refill_fetch_1_accessFault);
  assign MmuPlugin_logic_refill_onExit_BOOT = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_BOOT) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_BOOT));
  assign MmuPlugin_logic_refill_onExit_IDLE = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_IDLE) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_IDLE));
  assign MmuPlugin_logic_refill_onExit_CMD_0 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_CMD_0) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_CMD_0));
  assign MmuPlugin_logic_refill_onExit_CMD_1 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_CMD_1) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_CMD_1));
  assign MmuPlugin_logic_refill_onExit_RSP_0 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_RSP_0) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_RSP_0));
  assign MmuPlugin_logic_refill_onExit_RSP_1 = ((MmuPlugin_logic_refill_stateNext != MmuPlugin_logic_refill_RSP_1) && (MmuPlugin_logic_refill_stateReg == MmuPlugin_logic_refill_RSP_1));
  assign MmuPlugin_logic_refill_onEntry_BOOT = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_BOOT) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_BOOT));
  assign MmuPlugin_logic_refill_onEntry_IDLE = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_IDLE) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_IDLE));
  assign MmuPlugin_logic_refill_onEntry_CMD_0 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_CMD_0) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_CMD_0));
  assign MmuPlugin_logic_refill_onEntry_CMD_1 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_CMD_1) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_CMD_1));
  assign MmuPlugin_logic_refill_onEntry_RSP_0 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_RSP_0) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_RSP_0));
  assign MmuPlugin_logic_refill_onEntry_RSP_1 = ((MmuPlugin_logic_refill_stateNext == MmuPlugin_logic_refill_RSP_1) && (MmuPlugin_logic_refill_stateReg != MmuPlugin_logic_refill_RSP_1));
  always @(*) begin
    PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_stateReg;
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        if(PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_CSR_WRITE;
        end else begin
          if(PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
            PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_READ_LOW;
          end else begin
            if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
              PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_READ_LOW;
            end
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
        if(PerformanceCounterPlugin_logic_readPort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_CALC_LOW;
        end
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
        if(PerformanceCounterPlugin_logic_writePort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_IDLE;
          if(when_PerformanceCounterPlugin_l278) begin
            PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_READ_HIGH;
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
        if(PerformanceCounterPlugin_logic_readPort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_CALC_HIGH;
        end
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
        if(PerformanceCounterPlugin_logic_writePort_ready) begin
          PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_IDLE;
        end
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
        PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_IDLE;
      end
      default : begin
      end
    endcase
    if(PerformanceCounterPlugin_logic_fsm_wantStart) begin
      PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_IDLE;
    end
    if(PerformanceCounterPlugin_logic_fsm_wantKill) begin
      PerformanceCounterPlugin_logic_fsm_stateNext = PerformanceCounterPlugin_logic_fsm_BOOT;
    end
  end

  assign when_PerformanceCounterPlugin_l271 = PerformanceCounterPlugin_logic_fsm_counterReaded[7];
  assign when_PerformanceCounterPlugin_l278 = PerformanceCounterPlugin_logic_fsm_calc_sum[32];
  assign when_PerformanceCounterPlugin_l249 = (CsrAccessPlugin_bus_write_address[7] == 1'b0);
  assign when_PerformanceCounterPlugin_l255 = PerformanceCounterPlugin_logic_fsm_cmd_oh[1];
  assign PerformanceCounterPlugin_logic_fsm_onExit_BOOT = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_BOOT) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_BOOT));
  assign PerformanceCounterPlugin_logic_fsm_onExit_IDLE = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_IDLE) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_IDLE));
  assign PerformanceCounterPlugin_logic_fsm_onExit_READ_LOW = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_READ_LOW) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_READ_LOW));
  assign PerformanceCounterPlugin_logic_fsm_onExit_CALC_LOW = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_CALC_LOW) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_CALC_LOW));
  assign PerformanceCounterPlugin_logic_fsm_onExit_READ_HIGH = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_READ_HIGH) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_READ_HIGH));
  assign PerformanceCounterPlugin_logic_fsm_onExit_CALC_HIGH = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_CALC_HIGH) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_CALC_HIGH));
  assign PerformanceCounterPlugin_logic_fsm_onExit_CSR_WRITE = ((PerformanceCounterPlugin_logic_fsm_stateNext != PerformanceCounterPlugin_logic_fsm_CSR_WRITE) && (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_CSR_WRITE));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_BOOT = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_BOOT) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_BOOT));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_IDLE = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_IDLE) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_IDLE));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_READ_LOW = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_READ_LOW) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_READ_LOW));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_CALC_LOW = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_CALC_LOW) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_CALC_LOW));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_READ_HIGH = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_READ_HIGH) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_READ_HIGH));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_CALC_HIGH = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_CALC_HIGH) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_CALC_HIGH));
  assign PerformanceCounterPlugin_logic_fsm_onEntry_CSR_WRITE = ((PerformanceCounterPlugin_logic_fsm_stateNext == PerformanceCounterPlugin_logic_fsm_CSR_WRITE) && (PerformanceCounterPlugin_logic_fsm_stateReg != PerformanceCounterPlugin_logic_fsm_CSR_WRITE));
  assign PerformanceCounterPlugin_logic_fsm_done = (PerformanceCounterPlugin_logic_fsm_stateReg == PerformanceCounterPlugin_logic_fsm_IDLE);
  always @(*) begin
    CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_stateReg;
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        if(when_CsrAccessPlugin_l296) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_WRITE;
        end
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
        if(when_CsrAccessPlugin_l325) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_COMPLETION;
        end
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
        if(execute_ctrl2_down_isReady) begin
          CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_IDLE;
        end
      end
      default : begin
        if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
          if(when_CsrAccessPlugin_l212) begin
            CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_READ;
          end
          if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
            if(!CsrAccessPlugin_logic_fsm_inject_trapReg) begin
              CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_READ;
            end
          end
        end
      end
    endcase
    if(CsrAccessPlugin_logic_fsm_wantKill) begin
      CsrAccessPlugin_logic_fsm_stateNext = CsrAccessPlugin_logic_fsm_IDLE;
    end
  end

  assign when_CsrAccessPlugin_l296 = (! CsrAccessPlugin_bus_read_halt);
  assign when_CsrAccessPlugin_l325 = (! CsrAccessPlugin_bus_write_halt);
  assign when_CsrAccessPlugin_l212 = ((! CsrAccessPlugin_logic_fsm_inject_trap) && (! CsrAccessPlugin_bus_decode_trap));
  assign CsrAccessPlugin_logic_fsm_onExit_IDLE = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_IDLE) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_IDLE));
  assign CsrAccessPlugin_logic_fsm_onExit_READ = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_READ) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_READ));
  assign CsrAccessPlugin_logic_fsm_onExit_WRITE = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_WRITE) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_WRITE));
  assign CsrAccessPlugin_logic_fsm_onExit_COMPLETION = ((CsrAccessPlugin_logic_fsm_stateNext != CsrAccessPlugin_logic_fsm_COMPLETION) && (CsrAccessPlugin_logic_fsm_stateReg == CsrAccessPlugin_logic_fsm_COMPLETION));
  assign CsrAccessPlugin_logic_fsm_onEntry_IDLE = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_IDLE) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_IDLE));
  assign CsrAccessPlugin_logic_fsm_onEntry_READ = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_READ) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_READ));
  assign CsrAccessPlugin_logic_fsm_onEntry_WRITE = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_WRITE) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_WRITE));
  assign CsrAccessPlugin_logic_fsm_onEntry_COMPLETION = ((CsrAccessPlugin_logic_fsm_stateNext == CsrAccessPlugin_logic_fsm_COMPLETION) && (CsrAccessPlugin_logic_fsm_stateReg != CsrAccessPlugin_logic_fsm_COMPLETION));
  assign BtbPlugin_logic_ras_mem_stack_wr_en = (_zz_wr_en && 1'b1);
  assign BtbPlugin_logic_ras_mem_stack_wr_data = BtbPlugin_logic_ras_write_payload_data;
  assign LsuL1Plugin_logic_banks_0_mem_wr_en = (LsuL1Plugin_logic_banks_0_write_valid && 1'b1);
  assign LsuL1Plugin_logic_banks_0_mem_rd_en = (LsuL1Plugin_logic_banks_0_read_cmd_valid && 1'b1);
  assign LsuL1Plugin_logic_banks_1_mem_wr_en = (LsuL1Plugin_logic_banks_1_write_valid && 1'b1);
  assign LsuL1Plugin_logic_banks_1_mem_rd_en = (LsuL1Plugin_logic_banks_1_read_cmd_valid && 1'b1);
  assign LsuL1Plugin_logic_banks_2_mem_wr_en = (LsuL1Plugin_logic_banks_2_write_valid && 1'b1);
  assign LsuL1Plugin_logic_banks_2_mem_rd_en = (LsuL1Plugin_logic_banks_2_read_cmd_valid && 1'b1);
  assign LsuL1Plugin_logic_banks_3_mem_wr_en = (LsuL1Plugin_logic_banks_3_write_valid && 1'b1);
  assign LsuL1Plugin_logic_banks_3_mem_rd_en = (LsuL1Plugin_logic_banks_3_read_cmd_valid && 1'b1);
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_wr_en = (FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask[0] && 1'b1);
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_0_wr_data = {FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_wr_en = (FetchL1Plugin_logic_translationStorage_logic_sl_0_write_mask[1] && 1'b1);
  assign FetchL1Plugin_logic_translationStorage_logic_sl_0_ways_1_wr_data = {FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,FetchL1Plugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_wr_en = (FetchL1Plugin_logic_translationStorage_logic_sl_1_write_mask[0] && 1'b1);
  assign FetchL1Plugin_logic_translationStorage_logic_sl_1_ways_0_wr_data = {FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowUser,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowExecute,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowWrite,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_allowRead,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress,{FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress,FetchL1Plugin_logic_translationStorage_logic_sl_1_write_data_valid}}}}}};
  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_wr_en = (LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[0] && 1'b1);
  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_0_wr_data = {LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_wr_en = (LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[1] && 1'b1);
  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_1_wr_data = {LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_wr_en = (LsuPlugin_logic_translationStorage_logic_sl_0_write_mask[2] && 1'b1);
  assign LsuPlugin_logic_translationStorage_logic_sl_0_ways_2_wr_data = {LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_0_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_0_write_data_valid}}}}}};
  assign LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_wr_en = (LsuPlugin_logic_translationStorage_logic_sl_1_write_mask[0] && 1'b1);
  assign LsuPlugin_logic_translationStorage_logic_sl_1_ways_0_wr_data = {LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowUser,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowExecute,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowWrite,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_allowRead,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_physicalAddress,{LsuPlugin_logic_translationStorage_logic_sl_1_write_data_virtualAddress,LsuPlugin_logic_translationStorage_logic_sl_1_write_data_valid}}}}}};
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      MmuPlugin_logic_satp_mode <= 1'b0;
      MmuPlugin_logic_satp_ppn <= 20'h0;
      MmuPlugin_logic_status_mxr <= 1'b0;
      MmuPlugin_logic_status_sum <= 1'b0;
      CfuPlugin_logic_en <= 1'b0;
      CfuPlugin_logic_csr_stateId <= 3'b000;
      CfuPlugin_logic_csr_cfuIndex <= 4'b0000;
      CfuPlugin_logic_onFork_fired <= 1'b0;
      early0_DivPlugin_logic_processing_cmdSent <= 1'b0;
      early0_DivPlugin_logic_processing_unscheduleRequest <= 1'b0;
      FetchL1Plugin_logic_invalidate_counter <= 7'h0;
      FetchL1Plugin_logic_invalidate_firstEver <= 1'b1;
      FetchL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
      FetchL1Plugin_logic_refill_pushCounter <= 32'h0;
      FetchL1Plugin_logic_refill_onCmd_locked <= 1'b0;
      FetchL1Plugin_logic_refill_onRsp_wordIndex <= 3'b000;
      FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b1;
      FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid <= 1'b0;
      FetchL1Plugin_logic_ctrl_trapSent <= 1'b0;
      FetchL1Plugin_logic_ctrl_firstCycle <= 1'b1;
      FetchL1Plugin_logic_ctrl_onEvents_waiting <= 1'b0;
      PrivilegedPlugin_logic_harts_0_privilege <= 2'b11;
      PrivilegedPlugin_logic_harts_0_m_status_mie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_mpie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b00;
      PrivilegedPlugin_logic_harts_0_m_status_fs <= 2'b00;
      PrivilegedPlugin_logic_harts_0_m_status_tsr <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_tvm <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_tw <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_status_mprv <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_harts_0_m_ip_meip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ip_mtip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ip_msip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_meie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_mtie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ie_msie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_iam <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_bp <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_eu <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_es <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_ipf <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_lpf <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_edeleg_spf <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ideleg_st <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ideleg_se <= 1'b0;
      PrivilegedPlugin_logic_harts_0_m_ideleg_ss <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_cause_interrupt <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_cause_code <= 4'b0000;
      PrivilegedPlugin_logic_harts_0_s_status_sie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_status_spie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_status_spp <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ip_seipSoft <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ip_stip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ip_ssip <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ie_seie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ie_stie <= 1'b0;
      PrivilegedPlugin_logic_harts_0_s_ie_ssie <= 1'b0;
      BtbPlugin_logic_ras_ptr_push <= 2'b00;
      BtbPlugin_logic_ras_ptr_pop <= 2'b11;
      decode_ctrls_0_up_LANE_SEL_0_regNext <= 1'b0;
      PerformanceCounterPlugin_logic_ignoreNextCommit <= 1'b0;
      PerformanceCounterPlugin_logic_counters_cycle_value <= 8'h0;
      PerformanceCounterPlugin_logic_counters_cycle_mcounteren <= 1'b0;
      PerformanceCounterPlugin_logic_counters_cycle_scounteren <= 1'b0;
      PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit <= 1'b0;
      PerformanceCounterPlugin_logic_counters_instret_value <= 8'h0;
      PerformanceCounterPlugin_logic_counters_instret_mcounteren <= 1'b0;
      PerformanceCounterPlugin_logic_counters_instret_scounteren <= 1'b0;
      PerformanceCounterPlugin_logic_counters_instret_mcountinhibit <= 1'b0;
      _zz_PerformanceCounterPlugin_logic_counters_instret_value <= 1'b0;
      AlignerPlugin_logic_feeder_harts_0_dopId <= 10'h0;
      AlignerPlugin_logic_nobuffer_mask <= 1'b1;
      execute_ctrl3_up_CfuPlugin_logic_CFU_IN_FLIGHT_lane0 <= 1'b0;
      execute_ctrl4_up_CfuPlugin_logic_CFU_IN_FLIGHT_lane0 <= 1'b0;
      DecoderPlugin_logic_harts_0_uopId <= 16'h0;
      DecoderPlugin_logic_interrupt_buffered <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_0_regNext <= 1'b0;
      DispatchPlugin_logic_feeds_0_sent <= 1'b0;
      CsrRamPlugin_csrMapper_fired <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= 1'b0;
      execute_ctrl0_down_LANE_SEL_lane0_regNext <= 1'b0;
      execute_ctrl2_down_LANE_SEL_lane0_regNext <= 1'b0;
      BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      decode_ctrls_1_up_LANE_SEL_0 <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b1;
      LsuL1Plugin_logic_refill_pushCounter <= 32'h0;
      LsuL1Plugin_logic_refill_read_arbiter_lock <= 1'b0;
      LsuL1Plugin_logic_refill_read_wordIndex <= 3'b000;
      LsuL1Plugin_logic_refill_read_hadError <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b0;
      LsuL1Plugin_logic_writeback_read_arbiter_lock <= 1'b0;
      LsuL1Plugin_logic_writeback_read_wordIndex <= 3'b000;
      LsuL1Plugin_logic_writeback_read_slotReadLast_valid <= 1'b0;
      LsuL1Plugin_logic_writeback_write_arbiter_lock <= 1'b0;
      LsuL1Plugin_logic_writeback_write_wordIndex <= 3'b000;
      LsuL1Plugin_logic_writeback_write_bufferRead_rValid <= 1'b0;
      LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg <= 1'b0;
      LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg <= 1'b0;
      LsuL1Plugin_logic_lsu_rb1_onBanks_2_busyReg <= 1'b0;
      LsuL1Plugin_logic_lsu_rb1_onBanks_3_busyReg <= 1'b0;
      LsuL1Plugin_logic_lsu_ctrl_hazardReg <= 1'b0;
      LsuL1Plugin_logic_lsu_ctrl_flushHazardReg <= 1'b0;
      LsuL1Plugin_logic_initializer_counter <= 7'h0;
      TrapPlugin_logic_harts_0_interrupt_validBuffer <= 1'b0;
      TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated <= 1'b0;
      TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug <= 1'b0;
      LsuPlugin_logic_onAddress0_ls_storeId <= 12'h0;
      LsuPlugin_logic_onAddress0_access_waiter_valid <= 1'b0;
      execute_ctrl3_up_LsuL1_SEL_lane0 <= 1'b0;
      execute_ctrl4_up_LsuL1_SEL_lane0 <= 1'b0;
      LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b0;
      LsuPlugin_logic_onCtrl_io_allowIt <= 1'b0;
      LsuPlugin_logic_onCtrl_io_doItReg <= 1'b0;
      LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b0;
      LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b0;
      LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= 1'b0;
      LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b0;
      LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock <= 1'b0;
      LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat <= 3'b000;
      PcPlugin_logic_harts_0_self_id <= 10'h0;
      PcPlugin_logic_harts_0_self_increment <= 1'b0;
      PcPlugin_logic_harts_0_self_fault <= 1'b0;
      PcPlugin_logic_harts_0_self_state <= 32'h0;
      PcPlugin_logic_harts_0_holdReg <= 1'b1;
      HistoryPlugin_logic_onFetch_value <= 12'h0;
      FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value <= 1'b0;
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value <= 2'b00;
      MmuPlugin_logic_refill_cacheRefillAny <= 1'b0;
      MmuPlugin_logic_refill_load_rsp_valid <= 1'b0;
      MmuPlugin_logic_invalidate_busy <= 1'b0;
      PerformanceCounterPlugin_logic_interrupt_ip <= 1'b0;
      PerformanceCounterPlugin_logic_interrupt_ie <= 1'b0;
      PerformanceCounterPlugin_logic_interrupt_sup_deleg <= 1'b0;
      PerformanceCounterPlugin_logic_csrRead_fired <= 1'b0;
      PerformanceCounterPlugin_logic_csrWrite_fired <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b0;
      CsrAccessPlugin_logic_fsm_inject_sampled <= 1'b0;
      CsrRamPlugin_logic_readLogic_ohReg <= 3'b000;
      CsrRamPlugin_logic_readLogic_busy <= 1'b0;
      CsrRamPlugin_logic_flush_counter <= 5'h0;
      execute_ctrl1_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl2_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl3_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl4_up_LANE_SEL_lane0 <= 1'b0;
      execute_ctrl5_up_LANE_SEL_lane0 <= 1'b0;
      integer_RegFilePlugin_logic_initalizer_counter <= 6'h0;
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 <= 60'h0;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 <= 60'h0;
      fetch_logic_ctrls_1_up_valid <= 1'b0;
      fetch_logic_ctrls_2_up_valid <= 1'b0;
      decode_ctrls_1_up_valid <= 1'b0;
      LsuPlugin_logic_flusher_stateReg <= LsuPlugin_logic_flusher_IDLE;
      TrapPlugin_logic_harts_0_trap_fsm_stateReg <= TrapPlugin_logic_harts_0_trap_fsm_RESET;
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_BOOT;
      PerformanceCounterPlugin_logic_fsm_stateReg <= PerformanceCounterPlugin_logic_fsm_BOOT;
      CsrAccessPlugin_logic_fsm_stateReg <= CsrAccessPlugin_logic_fsm_IDLE;
    end else begin
      if(CfuPlugin_logic_bus_cmd_fire) begin
        CfuPlugin_logic_onFork_fired <= 1'b1;
      end
      if(when_CfuPlugin_l147) begin
        CfuPlugin_logic_onFork_fired <= 1'b0;
      end
      if(early0_DivPlugin_logic_processing_div_io_cmd_fire) begin
        early0_DivPlugin_logic_processing_cmdSent <= 1'b1;
      end
      if(execute_ctrl2_down_isReady) begin
        early0_DivPlugin_logic_processing_cmdSent <= 1'b0;
      end
      early0_DivPlugin_logic_processing_unscheduleRequest <= execute_lane0_ctrls_2_upIsCancel;
      if(execute_ctrl2_down_isReady) begin
        early0_DivPlugin_logic_processing_unscheduleRequest <= 1'b0;
      end
      if(FetchL1Plugin_logic_invalidate_done) begin
        FetchL1Plugin_logic_invalidate_firstEver <= 1'b0;
      end
      if(when_FetchL1Plugin_l204) begin
        FetchL1Plugin_logic_invalidate_counter <= FetchL1Plugin_logic_invalidate_counterIncr;
      end
      if(when_FetchL1Plugin_l211) begin
        FetchL1Plugin_logic_invalidate_counter <= 7'h0;
      end
      if(when_FetchL1Plugin_l255) begin
        if(_zz_when) begin
          FetchL1Plugin_logic_refill_slots_0_valid <= 1'b1;
          FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b0;
        end
        FetchL1Plugin_logic_refill_pushCounter <= (FetchL1Plugin_logic_refill_pushCounter + 32'h00000001);
      end
      if(FetchL1Plugin_logic_bus_cmd_valid) begin
        FetchL1Plugin_logic_refill_onCmd_locked <= 1'b1;
      end
      if(FetchL1Plugin_logic_bus_cmd_ready) begin
        FetchL1Plugin_logic_refill_onCmd_locked <= 1'b0;
      end
      if(FetchL1Plugin_logic_bus_cmd_ready) begin
        if(FetchL1Plugin_logic_refill_onCmd_oh[0]) begin
          FetchL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
        end
      end
      if(FetchL1Plugin_logic_bus_rsp_fire) begin
        FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b0;
      end
      if(FetchL1Plugin_logic_bus_rsp_valid) begin
        FetchL1Plugin_logic_refill_onRsp_wordIndex <= (FetchL1Plugin_logic_refill_onRsp_wordIndex + 3'b001);
        if(when_FetchL1Plugin_l330) begin
          FetchL1Plugin_logic_refill_onRsp_firstCycle <= 1'b1;
          FetchL1Plugin_logic_refill_slots_0_valid <= 1'b0;
        end
      end
      FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_valid <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_valid;
      if(FetchL1Plugin_logic_trapPort_valid) begin
        FetchL1Plugin_logic_ctrl_trapSent <= 1'b1;
      end
      if(fetch_logic_ctrls_2_up_isCancel) begin
        FetchL1Plugin_logic_ctrl_trapSent <= 1'b0;
      end
      if(fetch_logic_ctrls_2_up_isValid) begin
        FetchL1Plugin_logic_ctrl_firstCycle <= 1'b0;
      end
      if(when_FetchL1Plugin_l541) begin
        FetchL1Plugin_logic_ctrl_firstCycle <= 1'b1;
      end
      if(when_FetchL1Plugin_l549) begin
        FetchL1Plugin_logic_ctrl_onEvents_waiting <= 1'b0;
      end
      if(FetchL1Plugin_logic_events_miss) begin
        FetchL1Plugin_logic_ctrl_onEvents_waiting <= 1'b1;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((|FetchL1Plugin_logic_refill_slots_0_valid) && (! FetchL1Plugin_logic_invalidate_done)))); // FetchL1Plugin.scala:L556
        `else
          if(!(! ((|FetchL1Plugin_logic_refill_slots_0_valid) && (! FetchL1Plugin_logic_invalidate_done)))) begin
            $display("FAILURE "); // FetchL1Plugin.scala:L556
            $finish;
          end
        `endif
      `endif
      if(PrivilegedPlugin_logic_harts_0_xretAwayFromMachine) begin
        PrivilegedPlugin_logic_harts_0_m_status_mprv <= 1'b0;
      end
      PrivilegedPlugin_logic_harts_0_m_ip_meip <= PrivilegedPlugin_logic_harts_0_int_m_external;
      PrivilegedPlugin_logic_harts_0_m_ip_mtip <= PrivilegedPlugin_logic_harts_0_int_m_timer;
      PrivilegedPlugin_logic_harts_0_m_ip_msip <= PrivilegedPlugin_logic_harts_0_int_m_software;
      BtbPlugin_logic_ras_ptr_push <= (_zz_BtbPlugin_logic_ras_ptr_push - _zz_BtbPlugin_logic_ras_ptr_push_3);
      decode_ctrls_0_up_LANE_SEL_0_regNext <= decode_ctrls_0_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l50) begin
        decode_ctrls_0_up_LANE_SEL_0_regNext <= 1'b0;
      end
      if(when_PerformanceCounterPlugin_l45) begin
        PerformanceCounterPlugin_logic_ignoreNextCommit <= 1'b0;
      end
      PerformanceCounterPlugin_logic_counters_cycle_value <= (PerformanceCounterPlugin_logic_counters_cycle_value + _zz_PerformanceCounterPlugin_logic_counters_cycle_value);
      _zz_PerformanceCounterPlugin_logic_counters_instret_value <= ((! PerformanceCounterPlugin_logic_counters_instret_mcountinhibit) ? PerformanceCounterPlugin_logic_commitCount : 1'b0);
      PerformanceCounterPlugin_logic_counters_instret_value <= (PerformanceCounterPlugin_logic_counters_instret_value + _zz_PerformanceCounterPlugin_logic_counters_instret_value_1);
      if(when_AlignerPlugin_l171) begin
        AlignerPlugin_logic_feeder_harts_0_dopId <= (decode_ctrls_0_down_Decode_DOP_ID_0 + 10'h001);
      end
      if(when_AlignerPlugin_l292) begin
        AlignerPlugin_logic_nobuffer_mask <= AlignerPlugin_logic_nobuffer_remaningMask;
      end
      if(when_DecoderPlugin_l143) begin
        DecoderPlugin_logic_harts_0_uopId <= (DecoderPlugin_logic_harts_0_uopId + 16'h0001);
      end
      if(when_DecoderPlugin_l151) begin
        DecoderPlugin_logic_interrupt_buffered <= DecoderPlugin_logic_interrupt_async;
      end
      decode_ctrls_1_up_LANE_SEL_0_regNext <= decode_ctrls_1_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l50_1) begin
        decode_ctrls_1_up_LANE_SEL_0_regNext <= 1'b0;
      end
      if(DispatchPlugin_logic_feeds_0_sending) begin
        DispatchPlugin_logic_feeds_0_sent <= 1'b1;
      end
      if(decode_ctrls_1_up_isMoving) begin
        DispatchPlugin_logic_feeds_0_sent <= 1'b0;
      end
      if(when_CsrRamPlugin_l92) begin
        CsrRamPlugin_csrMapper_fired <= 1'b1;
      end
      if(CsrAccessPlugin_bus_write_moving) begin
        CsrRamPlugin_csrMapper_fired <= 1'b0;
      end
      decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= decode_ctrls_1_up_LANE_SEL_0;
      if(when_CtrlLaneApi_l50_2) begin
        decode_ctrls_1_up_LANE_SEL_0_regNext_1 <= 1'b0;
      end
      execute_ctrl0_down_LANE_SEL_lane0_regNext <= execute_ctrl0_down_LANE_SEL_lane0;
      if(when_CtrlLaneApi_l50_3) begin
        execute_ctrl0_down_LANE_SEL_lane0_regNext <= 1'b0;
      end
      execute_ctrl2_down_LANE_SEL_lane0_regNext <= execute_ctrl2_down_LANE_SEL_lane0;
      if(when_CtrlLaneApi_l50_4) begin
        execute_ctrl2_down_LANE_SEL_lane0_regNext <= 1'b0;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[0]))); // BtbPlugin.scala:L215
        `else
          if(!(! (fetch_logic_ctrls_1_up_isValid && fetch_logic_ctrls_1_down_BtbPlugin_logic_readCmd_HAZARDS[0]))) begin
            $display("FAILURE "); // BtbPlugin.scala:L215
            $finish;
          end
        `endif
      `endif
      if(fetch_logic_ctrls_1_up_isValid) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b1;
      end
      if(when_BtbPlugin_l233) begin
        BtbPlugin_logic_applyIt_correctionSent <= 1'b0;
      end
      if(when_AlignerPlugin_l298) begin
        AlignerPlugin_logic_nobuffer_mask <= 1'b1;
      end
      if(LsuL1Plugin_logic_refill_slots_0_loadedSet) begin
        LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b1;
      end
      if(LsuL1Plugin_logic_refill_slots_0_fire) begin
        LsuL1Plugin_logic_refill_slots_0_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_refill_push_valid) begin
        LsuL1Plugin_logic_refill_pushCounter <= (LsuL1Plugin_logic_refill_pushCounter + 32'h00000001);
      end
      if(when_LsuL1Plugin_l377) begin
        LsuL1Plugin_logic_refill_slots_0_valid <= 1'b1;
        LsuL1Plugin_logic_refill_slots_0_loaded <= 1'b0;
      end
      LsuL1Plugin_logic_refill_read_arbiter_lock <= LsuL1Plugin_logic_refill_read_arbiter_oh;
      if(LsuL1Plugin_logic_bus_read_cmd_fire) begin
        LsuL1Plugin_logic_refill_read_arbiter_lock <= 1'b0;
      end
      if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(LsuL1Plugin_logic_refill_read_writeReservation_win); // LsuL1Plugin.scala:L429
          `else
            if(!LsuL1Plugin_logic_refill_read_writeReservation_win) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L429
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l450) begin
        LsuL1Plugin_logic_refill_read_hadError <= 1'b1;
      end
      if(LsuL1Plugin_logic_bus_read_rsp_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(LsuL1Plugin_logic_refill_read_reservation_win); // LsuL1Plugin.scala:L459
          `else
            if(!LsuL1Plugin_logic_refill_read_reservation_win) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L459
              $finish;
            end
          `endif
        `endif
        if(LsuL1Plugin_logic_refill_read_rspWithData) begin
          LsuL1Plugin_logic_refill_read_wordIndex <= (LsuL1Plugin_logic_refill_read_wordIndex + 3'b001);
        end
        if(when_LsuL1Plugin_l463) begin
          LsuL1Plugin_logic_refill_read_hadError <= 1'b0;
        end
      end
      if(LsuL1Plugin_logic_writeback_slots_0_fire) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      end
      if(LsuL1Plugin_logic_writeback_slots_0_fire) begin
        LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b0;
      end
      if(when_LsuL1Plugin_l530) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b0;
      end
      if(when_LsuL1Plugin_l556) begin
        LsuL1Plugin_logic_writeback_slots_0_valid <= 1'b1;
        LsuL1Plugin_logic_writeback_slots_0_busy <= 1'b1;
      end
      LsuL1Plugin_logic_writeback_read_arbiter_lock <= LsuL1Plugin_logic_writeback_read_arbiter_oh;
      LsuL1Plugin_logic_writeback_read_wordIndex <= (LsuL1Plugin_logic_writeback_read_wordIndex + _zz_LsuL1Plugin_logic_writeback_read_wordIndex);
      if(when_LsuL1Plugin_l605) begin
        LsuL1Plugin_logic_writeback_read_arbiter_lock <= 1'b0;
      end
      LsuL1Plugin_logic_writeback_read_slotReadLast_valid <= LsuL1Plugin_logic_writeback_read_slotRead_valid;
      LsuL1Plugin_logic_writeback_write_arbiter_lock <= LsuL1Plugin_logic_writeback_write_arbiter_oh;
      LsuL1Plugin_logic_writeback_write_wordIndex <= (LsuL1Plugin_logic_writeback_write_wordIndex + _zz_LsuL1Plugin_logic_writeback_write_wordIndex);
      if(when_LsuL1Plugin_l676) begin
        LsuL1Plugin_logic_writeback_write_arbiter_lock <= 1'b0;
      end
      if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
        LsuL1Plugin_logic_writeback_write_bufferRead_rValid <= LsuL1Plugin_logic_writeback_write_bufferRead_valid;
      end
      if(LsuL1Plugin_logic_banks_0_usedByWriteback) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l735) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_0_busyReg <= 1'b0;
      end
      if(LsuL1Plugin_logic_banks_1_usedByWriteback) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l735_1) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_1_busyReg <= 1'b0;
      end
      if(LsuL1Plugin_logic_banks_2_usedByWriteback) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_2_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l735_2) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_2_busyReg <= 1'b0;
      end
      if(LsuL1Plugin_logic_banks_3_usedByWriteback) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_3_busyReg <= 1'b1;
      end
      if(when_LsuL1Plugin_l735_3) begin
        LsuL1Plugin_logic_lsu_rb1_onBanks_3_busyReg <= 1'b0;
      end
      LsuL1Plugin_logic_lsu_ctrl_hazardReg <= (execute_ctrl4_down_LsuL1_HAZARD_lane0 && execute_freeze_valid);
      LsuL1Plugin_logic_lsu_ctrl_flushHazardReg <= (execute_ctrl4_down_LsuL1_FLUSH_HAZARD_lane0 && execute_freeze_valid);
      if(execute_ctrl4_down_LsuL1_SEL_lane0) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((_zz_58 <= 3'b001)); // LsuL1Plugin.scala:L892
          `else
            if(!(_zz_58 <= 3'b001)) begin
              $display("FAILURE Multiple way hit ???"); // LsuL1Plugin.scala:L892
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l915) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((_zz_64 < 2'b10)); // LsuL1Plugin.scala:L916
          `else
            if(!(_zz_64 < 2'b10)) begin
              $display("FAILURE "); // LsuL1Plugin.scala:L916
              $finish;
            end
          `endif
        `endif
      end
      if(when_LsuL1Plugin_l1219) begin
        LsuL1Plugin_logic_initializer_counter <= (LsuL1Plugin_logic_initializer_counter + 7'h01);
      end
      TrapPlugin_logic_harts_0_interrupt_validBuffer <= TrapPlugin_logic_harts_0_interrupt_valid;
      if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidate_cmd_fire) begin
        TrapPlugin_logic_harts_0_trap_fsm_atsPorts_invalidated <= 1'b1;
      end
      LsuPlugin_logic_onAddress0_ls_storeId <= (LsuPlugin_logic_onAddress0_ls_storeId + _zz_LsuPlugin_logic_onAddress0_ls_storeId);
      if(when_LsuPlugin_l259) begin
        LsuPlugin_logic_onAddress0_access_waiter_valid <= 1'b0;
      end
      LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b1;
      if(execute_freeze_valid) begin
        LsuPlugin_logic_onCtrl_io_tooEarly <= 1'b0;
      end
      LsuPlugin_logic_onCtrl_io_allowIt <= 1'b0;
      if(when_LsuPlugin_l597) begin
        LsuPlugin_logic_onCtrl_io_allowIt <= 1'b1;
      end
      LsuPlugin_logic_onCtrl_io_doItReg <= LsuPlugin_logic_onCtrl_io_doIt;
      if(LsuPlugin_logic_bus_cmd_fire) begin
        LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b1;
      end
      if(when_LsuPlugin_l601) begin
        LsuPlugin_logic_onCtrl_io_cmdSent <= 1'b0;
      end
      if(LsuPlugin_logic_bus_rsp_toStream_valid) begin
        LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b1;
      end
      if(LsuPlugin_logic_onCtrl_io_rsp_fire) begin
        LsuPlugin_logic_bus_rsp_toStream_rValid <= 1'b0;
      end
      if(when_LsuPlugin_l685) begin
        if(execute_ctrl4_down_LsuL1_STORE_lane0) begin
          LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= 1'b0;
        end
      end
      if(when_LsuPlugin_l697) begin
        LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= 1'b0;
      end
      if(LsuPlugin_logic_onCtrl_rva_lrsc_capture) begin
        LsuPlugin_logic_onCtrl_rva_lrsc_reserved <= (! LsuPlugin_logic_onCtrl_rva_lrsc_reserved);
      end
      if(when_LsuPlugin_l938) begin
        if(when_LsuPlugin_l263) begin
          LsuPlugin_logic_onAddress0_access_waiter_valid <= 1'b1;
        end
      end
      if(when_LsuPlugin_l259_1) begin
        LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b0;
      end
      if(when_LsuPlugin_l945) begin
        if(when_LsuPlugin_l263_1) begin
          LsuPlugin_logic_onCtrl_hartRegulation_valid <= 1'b1;
        end
      end
      if(LsuL1TileLinkPlugin_logic_down_a_valid) begin
        LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock <= 1'b1;
      end
      if(LsuL1TileLinkPlugin_logic_down_a_fire) begin
        LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat <= (LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat + 3'b001);
        if(LsuL1TileLinkPlugin_logic_down_a_tracker_last) begin
          LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_beat <= 3'b000;
        end
      end
      if(when_LsuL1Bus_l151) begin
        LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_lock <= 1'b0;
      end
      PcPlugin_logic_harts_0_holdReg <= PcPlugin_logic_harts_0_holdComb;
      PcPlugin_logic_harts_0_self_state <= PcPlugin_logic_harts_0_output_payload_pc;
      PcPlugin_logic_harts_0_self_fault <= PcPlugin_logic_harts_0_output_payload_fault;
      PcPlugin_logic_harts_0_self_increment <= 1'b0;
      if(PcPlugin_logic_harts_0_output_fire) begin
        PcPlugin_logic_harts_0_self_increment <= 1'b1;
      end
      if(fetch_logic_ctrls_0_up_isFiring) begin
        PcPlugin_logic_harts_0_self_id <= (PcPlugin_logic_harts_0_self_id + 10'h001);
      end
      HistoryPlugin_logic_onFetch_value <= HistoryPlugin_logic_onFetch_valueNext;
      FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_value <= FetchL1Plugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
      LsuPlugin_logic_translationStorage_logic_sl_0_allocId_value <= LsuPlugin_logic_translationStorage_logic_sl_0_allocId_valueNext;
      MmuPlugin_logic_refill_cacheRefillAny <= ((MmuPlugin_logic_refill_cacheRefillAny || MmuPlugin_logic_refill_cacheRefillAnySet) && (! 1'b0));
      MmuPlugin_logic_refill_load_rsp_valid <= MmuPlugin_logic_accessBus_rsp_valid;
      if(when_MmuPlugin_l512) begin
        if(MmuPlugin_logic_invalidate_arbiter_io_output_valid) begin
          MmuPlugin_logic_invalidate_busy <= 1'b1;
        end
      end else begin
        if(when_MmuPlugin_l526) begin
          MmuPlugin_logic_invalidate_busy <= 1'b0;
        end
      end
      if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_fire) begin
        PerformanceCounterPlugin_logic_csrRead_fired <= 1'b1;
      end
      if(CsrAccessPlugin_bus_read_moving) begin
        PerformanceCounterPlugin_logic_csrRead_fired <= 1'b0;
      end
      if(PerformanceCounterPlugin_logic_fsm_csrWriteCmd_fire) begin
        PerformanceCounterPlugin_logic_csrWrite_fired <= 1'b1;
      end
      if(CsrAccessPlugin_bus_write_moving) begin
        PerformanceCounterPlugin_logic_csrWrite_fired <= 1'b0;
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && execute_lane0_ctrls_2_upIsCancel))); // CsrAccessPlugin.scala:L136
        `else
          if(!(! ((execute_ctrl2_up_LANE_SEL_lane0 && execute_ctrl2_down_CsrAccessPlugin_SEL_lane0) && execute_lane0_ctrls_2_upIsCancel))) begin
            $display("FAILURE CsrAccessPlugin saw forbidden select && cancel request"); // CsrAccessPlugin.scala:L136
            $finish;
          end
        `endif
      `endif
      CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b0;
      if(CsrAccessPlugin_logic_flushPort_valid) begin
        CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b1;
      end
      if(when_CsrAccessPlugin_l197) begin
        CsrAccessPlugin_logic_fsm_inject_flushReg <= 1'b0;
      end
      CsrAccessPlugin_logic_fsm_inject_sampled <= execute_freeze_valid;
      if(when_CsrAccessPlugin_l346) begin
        MmuPlugin_logic_status_mxr <= CsrAccessPlugin_bus_write_bits[19];
        MmuPlugin_logic_status_sum <= CsrAccessPlugin_bus_write_bits[18];
        PrivilegedPlugin_logic_harts_0_m_status_mpie <= CsrAccessPlugin_bus_write_bits[7];
        PrivilegedPlugin_logic_harts_0_m_status_mie <= CsrAccessPlugin_bus_write_bits[3];
        if(when_CsrService_l176) begin
          case(switch_PrivilegedPlugin_l549)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b11;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b01;
            end
            2'b00 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b00;
            end
            default : begin
            end
          endcase
        end
        PrivilegedPlugin_logic_harts_0_m_status_mprv <= CsrAccessPlugin_bus_write_bits[17];
        PrivilegedPlugin_logic_harts_0_m_status_fs <= CsrAccessPlugin_bus_write_bits[14 : 13];
        PrivilegedPlugin_logic_harts_0_m_status_tsr <= CsrAccessPlugin_bus_write_bits[22];
        PrivilegedPlugin_logic_harts_0_m_status_tvm <= CsrAccessPlugin_bus_write_bits[20];
        PrivilegedPlugin_logic_harts_0_m_status_tw <= CsrAccessPlugin_bus_write_bits[21];
        PrivilegedPlugin_logic_harts_0_s_status_spp <= CsrAccessPlugin_bus_write_bits[8 : 8];
        PrivilegedPlugin_logic_harts_0_s_status_spie <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_status_sie <= CsrAccessPlugin_bus_write_bits[1];
      end
      if(when_CsrAccessPlugin_l346_1) begin
        MmuPlugin_logic_status_mxr <= CsrAccessPlugin_bus_write_bits[19];
        MmuPlugin_logic_status_sum <= CsrAccessPlugin_bus_write_bits[18];
        PrivilegedPlugin_logic_harts_0_s_status_spp <= CsrAccessPlugin_bus_write_bits[8 : 8];
        PrivilegedPlugin_logic_harts_0_s_status_spie <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_status_sie <= CsrAccessPlugin_bus_write_bits[1];
        PrivilegedPlugin_logic_harts_0_m_status_fs <= CsrAccessPlugin_bus_write_bits[14 : 13];
      end
      if(when_CsrAccessPlugin_l353) begin
        if(when_CsrAccessPlugin_l346_2) begin
          MmuPlugin_logic_satp_mode <= CsrAccessPlugin_bus_write_bits[31 : 31];
          MmuPlugin_logic_satp_ppn <= CsrAccessPlugin_bus_write_bits[19 : 0];
        end
      end
      if(when_CsrAccessPlugin_l346_3) begin
        CfuPlugin_logic_en <= CsrAccessPlugin_bus_write_bits[31];
        CfuPlugin_logic_csr_stateId <= CsrAccessPlugin_bus_write_bits[18 : 16];
        CfuPlugin_logic_csr_cfuIndex <= CsrAccessPlugin_bus_write_bits[3 : 0];
      end
      if(when_CsrAccessPlugin_l346_4) begin
        PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= CsrAccessPlugin_bus_write_bits[31];
        PrivilegedPlugin_logic_harts_0_m_cause_code <= CsrAccessPlugin_bus_write_bits[3 : 0];
      end
      if(when_CsrAccessPlugin_l346_5) begin
        PrivilegedPlugin_logic_harts_0_s_ip_seipSoft <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_s_ip_stip <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_ip_ssip <= CsrAccessPlugin_bus_write_bits[1];
        PerformanceCounterPlugin_logic_interrupt_ip <= CsrAccessPlugin_bus_write_bits[13];
      end
      if(when_CsrAccessPlugin_l346_6) begin
        PrivilegedPlugin_logic_harts_0_m_ie_meie <= CsrAccessPlugin_bus_write_bits[11];
        PrivilegedPlugin_logic_harts_0_m_ie_mtie <= CsrAccessPlugin_bus_write_bits[7];
        PrivilegedPlugin_logic_harts_0_m_ie_msie <= CsrAccessPlugin_bus_write_bits[3];
        PrivilegedPlugin_logic_harts_0_s_ie_seie <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_s_ie_stie <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_s_ie_ssie <= CsrAccessPlugin_bus_write_bits[1];
        PerformanceCounterPlugin_logic_interrupt_ie <= CsrAccessPlugin_bus_write_bits[13];
      end
      if(when_CsrAccessPlugin_l346_7) begin
        PrivilegedPlugin_logic_harts_0_m_edeleg_iam <= CsrAccessPlugin_bus_write_bits[0];
        PrivilegedPlugin_logic_harts_0_m_edeleg_bp <= CsrAccessPlugin_bus_write_bits[3];
        PrivilegedPlugin_logic_harts_0_m_edeleg_eu <= CsrAccessPlugin_bus_write_bits[8];
        PrivilegedPlugin_logic_harts_0_m_edeleg_es <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_m_edeleg_ipf <= CsrAccessPlugin_bus_write_bits[12];
        PrivilegedPlugin_logic_harts_0_m_edeleg_lpf <= CsrAccessPlugin_bus_write_bits[13];
        PrivilegedPlugin_logic_harts_0_m_edeleg_spf <= CsrAccessPlugin_bus_write_bits[15];
      end
      if(when_CsrAccessPlugin_l346_8) begin
        PrivilegedPlugin_logic_harts_0_m_ideleg_se <= CsrAccessPlugin_bus_write_bits[9];
        PrivilegedPlugin_logic_harts_0_m_ideleg_st <= CsrAccessPlugin_bus_write_bits[5];
        PrivilegedPlugin_logic_harts_0_m_ideleg_ss <= CsrAccessPlugin_bus_write_bits[1];
        PerformanceCounterPlugin_logic_interrupt_sup_deleg <= CsrAccessPlugin_bus_write_bits[13];
      end
      if(when_CsrAccessPlugin_l346_9) begin
        PrivilegedPlugin_logic_harts_0_s_cause_interrupt <= CsrAccessPlugin_bus_write_bits[31];
        PrivilegedPlugin_logic_harts_0_s_cause_code <= CsrAccessPlugin_bus_write_bits[3 : 0];
      end
      if(when_CsrAccessPlugin_l346_10) begin
        if(when_CsrService_l176) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_se) begin
            PrivilegedPlugin_logic_harts_0_s_ie_seie <= CsrAccessPlugin_bus_write_bits[9];
          end
        end
        if(when_CsrService_l176) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_st) begin
            PrivilegedPlugin_logic_harts_0_s_ie_stie <= CsrAccessPlugin_bus_write_bits[5];
          end
        end
        if(when_CsrService_l176) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_ss) begin
            PrivilegedPlugin_logic_harts_0_s_ie_ssie <= CsrAccessPlugin_bus_write_bits[1];
          end
        end
      end
      if(when_CsrAccessPlugin_l346_11) begin
        if(when_CsrService_l176) begin
          if(PrivilegedPlugin_logic_harts_0_m_ideleg_ss) begin
            PrivilegedPlugin_logic_harts_0_s_ip_ssip <= CsrAccessPlugin_bus_write_bits[1];
          end
        end
      end
      if(when_CsrAccessPlugin_l346_12) begin
        PerformanceCounterPlugin_logic_counters_cycle_mcounteren <= CsrAccessPlugin_bus_write_bits[0];
        PerformanceCounterPlugin_logic_counters_instret_mcounteren <= CsrAccessPlugin_bus_write_bits[2];
      end
      if(when_CsrAccessPlugin_l346_13) begin
        PerformanceCounterPlugin_logic_counters_cycle_scounteren <= CsrAccessPlugin_bus_write_bits[0];
        PerformanceCounterPlugin_logic_counters_instret_scounteren <= CsrAccessPlugin_bus_write_bits[2];
      end
      if(when_CsrAccessPlugin_l346_14) begin
        PerformanceCounterPlugin_logic_counters_cycle_mcountinhibit <= CsrAccessPlugin_bus_write_bits[0];
        PerformanceCounterPlugin_logic_counters_instret_mcountinhibit <= CsrAccessPlugin_bus_write_bits[2];
      end
      CsrRamPlugin_logic_readLogic_ohReg <= (CsrRamPlugin_logic_readLogic_port_cmd_valid ? CsrRamPlugin_logic_readLogic_oh : 3'b000);
      CsrRamPlugin_logic_readLogic_busy <= CsrRamPlugin_logic_readLogic_port_cmd_valid;
      CsrRamPlugin_logic_flush_counter <= (CsrRamPlugin_logic_flush_counter + _zz_CsrRamPlugin_logic_flush_counter);
      if(when_RegFilePlugin_l130) begin
        integer_RegFilePlugin_logic_initalizer_counter <= (integer_RegFilePlugin_logic_initalizer_counter + 6'h01);
      end
      _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_2 <= _zz_WhiteboxerPlugin_logic_perf_executeFreezedCounter_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchHazardsCounter_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_0_1;
      _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_2 <= _zz_WhiteboxerPlugin_logic_perf_candidatesCountCounters_1_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_0_1;
      _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_2 <= _zz_WhiteboxerPlugin_logic_perf_dispatchFeedCounters_1_1;
      if(fetch_logic_ctrls_1_up_forgetOne) begin
        fetch_logic_ctrls_1_up_valid <= 1'b0;
      end
      if(fetch_logic_ctrls_0_down_isReady) begin
        fetch_logic_ctrls_1_up_valid <= fetch_logic_ctrls_0_down_isValid;
      end
      if(fetch_logic_ctrls_2_up_forgetOne) begin
        fetch_logic_ctrls_2_up_valid <= 1'b0;
      end
      if(fetch_logic_ctrls_1_down_isReady) begin
        fetch_logic_ctrls_2_up_valid <= fetch_logic_ctrls_1_down_isValid;
      end
      if(decode_ctrls_0_down_isReady) begin
        decode_ctrls_1_up_valid <= decode_ctrls_0_down_isValid;
      end
      if(decode_ctrls_0_down_isReady) begin
        decode_ctrls_1_up_LANE_SEL_0 <= decode_ctrls_0_down_LANE_SEL_0;
      end
      if(when_DecodePipelinePlugin_l70) begin
        decode_ctrls_1_up_LANE_SEL_0 <= 1'b0;
      end
      if(execute_ctrl0_down_isReady) begin
        execute_ctrl1_up_LANE_SEL_lane0 <= execute_ctrl0_down_LANE_SEL_lane0;
      end
      if(execute_ctrl1_down_isReady) begin
        execute_ctrl2_up_LANE_SEL_lane0 <= execute_ctrl1_down_LANE_SEL_lane0;
      end
      if(execute_ctrl2_down_isReady) begin
        execute_ctrl3_up_LANE_SEL_lane0 <= execute_ctrl2_down_LANE_SEL_lane0;
        execute_ctrl3_up_CfuPlugin_logic_CFU_IN_FLIGHT_lane0 <= execute_ctrl2_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0;
        execute_ctrl3_up_LsuL1_SEL_lane0 <= execute_ctrl2_down_LsuL1_SEL_lane0;
      end
      if(execute_ctrl3_down_isReady) begin
        execute_ctrl4_up_LANE_SEL_lane0 <= execute_ctrl3_down_LANE_SEL_lane0;
        execute_ctrl4_up_CfuPlugin_logic_CFU_IN_FLIGHT_lane0 <= execute_ctrl3_down_CfuPlugin_logic_CFU_IN_FLIGHT_lane0;
        execute_ctrl4_up_LsuL1_SEL_lane0 <= execute_ctrl3_down_LsuL1_SEL_lane0;
      end
      if(execute_ctrl4_down_isReady) begin
        execute_ctrl5_up_LANE_SEL_lane0 <= execute_ctrl4_down_LANE_SEL_lane0;
      end
      LsuPlugin_logic_flusher_stateReg <= LsuPlugin_logic_flusher_stateNext;
      TrapPlugin_logic_harts_0_trap_fsm_stateReg <= TrapPlugin_logic_harts_0_trap_fsm_stateNext;
      case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
        TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
          TrapPlugin_logic_harts_0_trap_fsm_trapEnterDebug <= 1'b0;
          if(!when_TrapPlugin_l409) begin
            case(TrapPlugin_logic_harts_0_trap_pending_state_code)
              4'b0000 : begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert((! TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid)); // TrapPlugin.scala:L431
                  `else
                    if(!(! TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid)) begin
                      $display("FAILURE "); // TrapPlugin.scala:L431
                      $finish;
                    end
                  `endif
                `endif
              end
              4'b0001 : begin
              end
              4'b0010 : begin
              end
              4'b0100 : begin
              end
              4'b0101 : begin
              end
              4'b1000 : begin
              end
              4'b0110 : begin
              end
              4'b0111 : begin
              end
              default : begin
                `ifndef SYNTHESIS
                  `ifdef FORMAL
                    assert(1'b0); // TrapPlugin.scala:L482
                  `else
                    if(!1'b0) begin
                      $display("FAILURE Unexpected trap reason"); // TrapPlugin.scala:L482
                      $finish;
                    end
                  `endif
                `endif
              end
            endcase
          end
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
          PrivilegedPlugin_logic_harts_0_privilege <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege;
          case(TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_targetPrivilege)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mie <= 1'b0;
              PrivilegedPlugin_logic_harts_0_m_status_mpie <= PrivilegedPlugin_logic_harts_0_m_status_mie;
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= PrivilegedPlugin_logic_harts_0_privilege;
              PrivilegedPlugin_logic_harts_0_m_cause_code <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
              PrivilegedPlugin_logic_harts_0_m_cause_interrupt <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_harts_0_s_status_sie <= 1'b0;
              PrivilegedPlugin_logic_harts_0_s_status_spie <= PrivilegedPlugin_logic_harts_0_s_status_sie;
              PrivilegedPlugin_logic_harts_0_s_status_spp <= PrivilegedPlugin_logic_harts_0_privilege[0 : 0];
              PrivilegedPlugin_logic_harts_0_s_cause_code <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_code;
              PrivilegedPlugin_logic_harts_0_s_cause_interrupt <= TrapPlugin_logic_harts_0_trap_fsm_buffer_trap_interrupt;
            end
            default : begin
            end
          endcase
        end
        TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
          PrivilegedPlugin_logic_harts_0_privilege <= TrapPlugin_logic_harts_0_trap_pending_xret_targetPrivilege;
          case(switch_TrapPlugin_l655)
            2'b11 : begin
              PrivilegedPlugin_logic_harts_0_m_status_mpp <= 2'b00;
              PrivilegedPlugin_logic_harts_0_m_status_mie <= PrivilegedPlugin_logic_harts_0_m_status_mpie;
              PrivilegedPlugin_logic_harts_0_m_status_mpie <= 1'b1;
            end
            2'b01 : begin
              PrivilegedPlugin_logic_harts_0_s_status_spp <= 1'b0;
              PrivilegedPlugin_logic_harts_0_s_status_sie <= PrivilegedPlugin_logic_harts_0_s_status_spie;
              PrivilegedPlugin_logic_harts_0_s_status_spie <= 1'b1;
            end
            default : begin
            end
          endcase
        end
        TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
        end
        TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
        end
        default : begin
        end
      endcase
      MmuPlugin_logic_refill_stateReg <= MmuPlugin_logic_refill_stateNext;
      PerformanceCounterPlugin_logic_fsm_stateReg <= PerformanceCounterPlugin_logic_fsm_stateNext;
      case(PerformanceCounterPlugin_logic_fsm_stateReg)
        PerformanceCounterPlugin_logic_fsm_IDLE : begin
        end
        PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
        end
        PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
          if(when_PerformanceCounterPlugin_l271) begin
            if(_zz_PerformanceCounterPlugin_logic_fsm_cmd_address) begin
              PerformanceCounterPlugin_logic_counters_cycle_value[7] <= 1'b0;
            end
            if(_zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1) begin
              PerformanceCounterPlugin_logic_counters_instret_value[7] <= 1'b0;
            end
          end
        end
        PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
        end
        PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
        end
        PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
          if(when_PerformanceCounterPlugin_l249) begin
            if(_zz_PerformanceCounterPlugin_logic_fsm_cmd_address) begin
              PerformanceCounterPlugin_logic_counters_cycle_value <= _zz_PerformanceCounterPlugin_logic_counters_cycle_value_2[7:0];
              PerformanceCounterPlugin_logic_counters_cycle_value[7] <= 1'b0;
            end
            if(_zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1) begin
              PerformanceCounterPlugin_logic_counters_instret_value <= _zz_PerformanceCounterPlugin_logic_counters_instret_value_2[7:0];
              PerformanceCounterPlugin_logic_counters_instret_value[7] <= 1'b0;
            end
          end
          if(when_PerformanceCounterPlugin_l255) begin
            PerformanceCounterPlugin_logic_ignoreNextCommit <= 1'b1;
          end
        end
        default : begin
        end
      endcase
      CsrAccessPlugin_logic_fsm_stateReg <= CsrAccessPlugin_logic_fsm_stateNext;
      case(CsrAccessPlugin_logic_fsm_stateReg)
        CsrAccessPlugin_logic_fsm_READ : begin
        end
        CsrAccessPlugin_logic_fsm_WRITE : begin
        end
        CsrAccessPlugin_logic_fsm_COMPLETION : begin
        end
        default : begin
          if(CsrAccessPlugin_logic_fsm_inject_onDecodeDo) begin
            if(CsrAccessPlugin_logic_fsm_inject_sampled) begin
              if(CsrAccessPlugin_logic_fsm_inject_trapReg) begin
                CsrAccessPlugin_logic_fsm_inject_unfreeze <= execute_freeze_valid;
              end
            end
          end
        end
      endcase
      case(CsrAccessPlugin_logic_fsm_stateNext)
        CsrAccessPlugin_logic_fsm_READ : begin
        end
        CsrAccessPlugin_logic_fsm_WRITE : begin
        end
        CsrAccessPlugin_logic_fsm_COMPLETION : begin
          CsrAccessPlugin_logic_fsm_inject_unfreeze <= 1'b1;
        end
        default : begin
        end
      endcase
      BtbPlugin_logic_ras_ptr_pop <= BtbPlugin_logic_ras_ptr_pop_aheadValue;
    end
  end

  always @(posedge litex_clk) begin
    early0_DivPlugin_logic_processing_divRevertResult <= ((execute_ctrl2_down_RsUnsignedPlugin_RS1_REVERT_lane0 ^ (execute_ctrl2_down_RsUnsignedPlugin_RS2_REVERT_lane0 && (! execute_ctrl2_down_DivPlugin_REM_lane0))) && (! (((execute_ctrl2_down_RsUnsignedPlugin_RS2_FORMATED_lane0 == 32'h0) && execute_ctrl2_down_RsUnsignedPlugin_RS2_SIGNED_lane0) && (! execute_ctrl2_down_DivPlugin_REM_lane0))));
    if(when_FetchL1Plugin_l255) begin
      if(_zz_when) begin
        FetchL1Plugin_logic_refill_slots_0_address <= FetchL1Plugin_logic_refill_start_address;
        FetchL1Plugin_logic_refill_slots_0_isIo <= FetchL1Plugin_logic_refill_start_isIo;
        FetchL1Plugin_logic_refill_slots_0_wayToAllocate <= FetchL1Plugin_logic_refill_start_wayToAllocate;
        FetchL1Plugin_logic_refill_slots_0_priority <= FetchL1Plugin_logic_refill_slots_0_valid;
      end
    end
    if(when_FetchL1Plugin_l276) begin
      FetchL1Plugin_logic_refill_onCmd_lockedOh <= FetchL1Plugin_logic_refill_onCmd_propoedOh;
    end
    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_address <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_address;
    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_0 <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_0;
    FetchL1Plugin_logic_ctrl_plruLogic_buffer_regNext_payload_data_1 <= FetchL1Plugin_logic_ctrl_plruLogic_buffer_payload_data_1;
    PrivilegedPlugin_logic_harts_0_s_ip_seipInput <= PrivilegedPlugin_logic_harts_0_int_s_external;
    if(BtbPlugin_logic_ras_readIt) begin
      BtbPlugin_logic_ras_read <= BtbPlugin_logic_ras_mem_stack_rd_data;
    end
    LsuL1Plugin_logic_refill_slots_0_loadedCounter <= (LsuL1Plugin_logic_refill_slots_0_loadedCounter + ((LsuL1Plugin_logic_refill_slots_0_loaded && (! LsuL1Plugin_logic_refill_slots_0_loadedDone)) && (! execute_freeze_valid)));
    if(when_LsuL1Plugin_l381) begin
      LsuL1Plugin_logic_refill_slots_0_address <= LsuL1Plugin_logic_refill_push_payload_address;
      LsuL1Plugin_logic_refill_slots_0_way <= LsuL1Plugin_logic_refill_push_payload_way;
      LsuL1Plugin_logic_refill_slots_0_cmdSent <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_loadedCounter <= 1'b0;
      LsuL1Plugin_logic_refill_slots_0_victim <= LsuL1Plugin_logic_refill_push_payload_victim;
      LsuL1Plugin_logic_refill_slots_0_dirty <= LsuL1Plugin_logic_refill_push_payload_dirty;
    end
    if(LsuL1Plugin_logic_refill_read_arbiter_oh[0]) begin
      if(LsuL1Plugin_logic_bus_read_cmd_ready) begin
        LsuL1Plugin_logic_refill_slots_0_cmdSent <= 1'b1;
      end
    end
    LsuL1Plugin_logic_writeback_slots_0_timer_counter <= (LsuL1Plugin_logic_writeback_slots_0_timer_counter + ((! LsuL1Plugin_logic_writeback_slots_0_timer_done) && (! execute_freeze_valid)));
    if(when_LsuL1Plugin_l561) begin
      LsuL1Plugin_logic_writeback_slots_0_address <= LsuL1Plugin_logic_writeback_push_payload_address;
      LsuL1Plugin_logic_writeback_slots_0_way <= LsuL1Plugin_logic_writeback_push_payload_way;
      LsuL1Plugin_logic_writeback_slots_0_timer_counter <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_writeCmdDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_readCmdDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_readRspDone <= 1'b0;
      LsuL1Plugin_logic_writeback_slots_0_victimBufferReady <= 1'b0;
    end
    if(when_LsuL1Plugin_l605) begin
      if(LsuL1Plugin_logic_writeback_read_arbiter_oh[0]) begin
        LsuL1Plugin_logic_writeback_slots_0_readCmdDone <= 1'b1;
      end
    end
    if(LsuL1Plugin_logic_writeback_read_slotRead_valid) begin
      LsuL1Plugin_logic_refill_slots_0_victim[0] <= 1'b0;
    end
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last <= LsuL1Plugin_logic_writeback_read_slotRead_payload_last;
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_wordIndex <= LsuL1Plugin_logic_writeback_read_slotRead_payload_wordIndex;
    LsuL1Plugin_logic_writeback_read_slotReadLast_payload_way <= LsuL1Plugin_logic_writeback_read_slotRead_payload_way;
    if(LsuL1Plugin_logic_writeback_read_slotReadLast_valid) begin
      LsuL1Plugin_logic_writeback_slots_0_victimBufferReady <= 1'b1;
      if(LsuL1Plugin_logic_writeback_read_slotReadLast_payload_last) begin
        LsuL1Plugin_logic_writeback_slots_0_readRspDone <= 1'b1;
      end
    end
    if(when_LsuL1Plugin_l676) begin
      if(LsuL1Plugin_logic_writeback_write_arbiter_oh[0]) begin
        LsuL1Plugin_logic_writeback_slots_0_writeCmdDone <= 1'b1;
      end
    end
    if(LsuL1Plugin_logic_writeback_write_bufferRead_ready) begin
      LsuL1Plugin_logic_writeback_write_bufferRead_rData_address <= LsuL1Plugin_logic_writeback_write_bufferRead_payload_address;
      LsuL1Plugin_logic_writeback_write_bufferRead_rData_last <= LsuL1Plugin_logic_writeback_write_bufferRead_payload_last;
    end
    if(TrapPlugin_logic_harts_0_trap_pending_arbiter_down_valid) begin
      TrapPlugin_logic_harts_0_trap_pending_state_exception <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_exception;
      TrapPlugin_logic_harts_0_trap_pending_state_tval <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_tval;
      TrapPlugin_logic_harts_0_trap_pending_state_code <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_code;
      TrapPlugin_logic_harts_0_trap_pending_state_arg <= TrapPlugin_logic_harts_0_trap_pending_arbiter_down_payload_arg;
    end
    if(TrapPlugin_logic_harts_0_trap_trigger_valid) begin
      TrapPlugin_logic_harts_0_trap_pending_pc <= execute_ctrl4_down_PC_lane0;
      TrapPlugin_logic_harts_0_trap_pending_history <= execute_ctrl4_down_Prediction_BRANCH_HISTORY_lane0;
      TrapPlugin_logic_harts_0_trap_pending_slices <= (1'b0 + 1'b1);
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_valid <= TrapPlugin_logic_harts_0_interrupt_valid;
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_code <= TrapPlugin_logic_harts_0_interrupt_code;
    end
    if(TrapPlugin_logic_harts_0_trap_fsm_buffer_sampleIt) begin
      TrapPlugin_logic_harts_0_trap_fsm_buffer_i_targetPrivilege <= TrapPlugin_logic_harts_0_interrupt_targetPrivilege;
    end
    TrapPlugin_logic_harts_0_trap_fsm_jumpTarget <= (TrapPlugin_logic_harts_0_trap_pending_pc + _zz_TrapPlugin_logic_harts_0_trap_fsm_jumpTarget);
    if(when_TrapPlugin_l556) begin
      TrapPlugin_logic_harts_0_trap_fsm_readed <= TrapPlugin_logic_harts_0_crsPorts_read_data;
    end
    if(LsuPlugin_logic_onAddress0_flush_port_fire) begin
      LsuPlugin_logic_flusher_cmdCounter <= (LsuPlugin_logic_flusher_cmdCounter + 7'h01);
    end
    if(LsuPlugin_logic_bus_rsp_toStream_ready) begin
      LsuPlugin_logic_bus_rsp_toStream_rData_error <= LsuPlugin_logic_bus_rsp_toStream_payload_error;
      LsuPlugin_logic_bus_rsp_toStream_rData_data <= LsuPlugin_logic_bus_rsp_toStream_payload_data;
    end
    LsuPlugin_logic_onCtrl_rva_srcBuffer <= execute_ctrl4_down_LsuPlugin_logic_onCtrl_loadData_RESULT_lane0;
    LsuPlugin_logic_onCtrl_rva_aluBuffer <= LsuPlugin_logic_onCtrl_rva_alu_result;
    _zz_LsuPlugin_logic_onCtrl_rva_delay_0 <= (! execute_freeze_valid);
    _zz_LsuPlugin_logic_onCtrl_rva_delay_1 <= _zz_LsuPlugin_logic_onCtrl_rva_delay_0;
    if(!when_LsuPlugin_l697) begin
      LsuPlugin_logic_onCtrl_rva_lrsc_age <= (LsuPlugin_logic_onCtrl_rva_lrsc_age + _zz_LsuPlugin_logic_onCtrl_rva_lrsc_age);
    end
    if(LsuPlugin_logic_onCtrl_rva_lrsc_capture) begin
      LsuPlugin_logic_onCtrl_rva_lrsc_address <= execute_ctrl4_down_LsuL1_PHYSICAL_ADDRESS_lane0;
      LsuPlugin_logic_onCtrl_rva_lrsc_age <= 6'h0;
    end
    if(when_LsuPlugin_l901) begin
      LsuPlugin_logic_flusher_cmdCounter <= {1'd0, _zz_LsuPlugin_logic_flusher_cmdCounter};
    end
    if(when_LsuPlugin_l938) begin
      if(when_LsuPlugin_l263) begin
        LsuPlugin_logic_onAddress0_access_waiter_refill <= execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
      end
    end
    if(when_LsuPlugin_l945) begin
      if(when_LsuPlugin_l263_1) begin
        LsuPlugin_logic_onCtrl_hartRegulation_refill <= execute_ctrl4_down_LsuL1_WAIT_REFILL_lane0;
      end
    end
    LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_selReg <= LsuL1Plugin_logic_bus_toTilelink_nonCoherent_onA_sel;
    MmuPlugin_logic_refill_load_rsp_payload_data <= MmuPlugin_logic_accessBus_rsp_payload_data;
    MmuPlugin_logic_refill_load_rsp_payload_error <= MmuPlugin_logic_accessBus_rsp_payload_error;
    MmuPlugin_logic_refill_load_rsp_payload_redo <= MmuPlugin_logic_accessBus_rsp_payload_redo;
    MmuPlugin_logic_refill_load_rsp_payload_waitAny <= MmuPlugin_logic_accessBus_rsp_payload_waitAny;
    if(when_MmuPlugin_l512) begin
      MmuPlugin_logic_invalidate_counter <= 5'h0;
    end else begin
      MmuPlugin_logic_invalidate_counter <= (MmuPlugin_logic_invalidate_counter + 5'h01);
    end
    _zz_PerformanceCounterPlugin_logic_events_sums_0 <= early0_BranchPlugin_logic_events_branchMiss;
    _zz_PerformanceCounterPlugin_logic_events_sums_1 <= early0_BranchPlugin_logic_events_branchCount;
    _zz_PerformanceCounterPlugin_logic_events_sums_2 <= LsuPlugin_logic_events_waiting;
    _zz_PerformanceCounterPlugin_logic_events_sums_3 <= LsuL1Plugin_logic_events_loadAccess;
    _zz_PerformanceCounterPlugin_logic_events_sums_4 <= LsuL1Plugin_logic_events_loadMiss;
    _zz_PerformanceCounterPlugin_logic_events_sums_5 <= FetchL1Plugin_logic_events_access;
    _zz_PerformanceCounterPlugin_logic_events_sums_6 <= FetchL1Plugin_logic_events_miss;
    _zz_PerformanceCounterPlugin_logic_events_sums_7 <= FetchL1Plugin_logic_events_waiting;
    _zz_PerformanceCounterPlugin_logic_events_sums_8 <= PerformanceCounterPlugin_logic_eventCycles;
    _zz_PerformanceCounterPlugin_logic_events_sums_9 <= PerformanceCounterPlugin_logic_eventInstructions_0;
    _zz_PerformanceCounterPlugin_logic_events_sums_10 <= DispatchPlugin_logic_events_frontendStall;
    _zz_PerformanceCounterPlugin_logic_events_sums_11 <= DispatchPlugin_logic_events_backendStall;
    _zz_PerformanceCounterPlugin_logic_events_sums_12 <= MmuPlugin_logic_refill_events_onStorage_0_waiting;
    _zz_PerformanceCounterPlugin_logic_events_sums_13 <= MmuPlugin_logic_refill_events_onStorage_1_waiting;
    CsrAccessPlugin_logic_fsm_interface_read <= ((execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 && (! CsrAccessPlugin_logic_fsm_inject_trap)) && CsrAccessPlugin_logic_fsm_inject_csrRead);
    CsrAccessPlugin_logic_fsm_interface_write <= ((execute_ctrl2_down_CsrAccessPlugin_SEL_lane0 && (! CsrAccessPlugin_logic_fsm_inject_trap)) && CsrAccessPlugin_logic_fsm_inject_csrWrite);
    CsrAccessPlugin_logic_fsm_inject_trapReg <= CsrAccessPlugin_logic_fsm_inject_trap;
    CsrAccessPlugin_logic_fsm_inject_busTrapReg <= CsrAccessPlugin_bus_decode_trap;
    CsrAccessPlugin_logic_fsm_inject_busTrapCodeReg <= CsrAccessPlugin_bus_decode_trapCode;
    CsrAccessPlugin_logic_fsm_interface_onWriteBits <= CsrAccessPlugin_logic_fsm_writeLogic_alu_result;
    if(fetch_logic_ctrls_0_down_isReady) begin
      fetch_logic_ctrls_1_up_Fetch_WORD_PC <= fetch_logic_ctrls_0_down_Fetch_WORD_PC;
      fetch_logic_ctrls_1_up_Fetch_PC_FAULT <= fetch_logic_ctrls_0_down_Fetch_PC_FAULT;
      fetch_logic_ctrls_1_up_Fetch_ID <= fetch_logic_ctrls_0_down_Fetch_ID;
      _zz_1 <= 1'b0;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_VALID;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0 <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_0;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_1 <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_PLRU_BYPASS_DATA_1;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE;
      fetch_logic_ctrls_1_up_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS <= fetch_logic_ctrls_0_down_FetchL1Plugin_logic_cmd_TAGS_UPDATE_ADDRESS;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_HASH <= fetch_logic_ctrls_0_down_GSharePlugin_logic_HASH;
      fetch_logic_ctrls_1_up_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_0_down_Prediction_BRANCH_HISTORY;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_valid <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_valid;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_address <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_address;
      fetch_logic_ctrls_1_up_GSharePlugin_logic_BYPASS_payload_data_0 <= fetch_logic_ctrls_0_down_GSharePlugin_logic_BYPASS_payload_data_0;
      fetch_logic_ctrls_1_up_BtbPlugin_logic_readCmd_HAZARDS <= fetch_logic_ctrls_0_down_BtbPlugin_logic_readCmd_HAZARDS;
    end
    if(fetch_logic_ctrls_1_down_isReady) begin
      fetch_logic_ctrls_2_up_Fetch_WORD_PC <= fetch_logic_ctrls_1_down_Fetch_WORD_PC;
      fetch_logic_ctrls_2_up_Fetch_PC_FAULT <= fetch_logic_ctrls_1_down_Fetch_PC_FAULT;
      fetch_logic_ctrls_2_up_Fetch_ID <= fetch_logic_ctrls_1_down_Fetch_ID;
      fetch_logic_ctrls_2_up_Prediction_BRANCH_HISTORY <= fetch_logic_ctrls_1_down_Prediction_BRANCH_HISTORY;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_0_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_0_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_1_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_1_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_2_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_2_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_2_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_2_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_3_loaded <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_loaded;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_3_error <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_error;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_TAGS_3_address <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_TAGS_3_address;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_PLRU_BYPASSED_1 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_PLRU_BYPASSED_1;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_1 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_1;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_2 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_2;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_BANKS_MUXES_3 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_BANKS_MUXES_3;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_HAZARD <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_HAZARD;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_0 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_0;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_1 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_1;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_2 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_2;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HITS_3 <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HITS_3;
      fetch_logic_ctrls_2_up_MMU_BYPASS_TRANSLATION <= fetch_logic_ctrls_1_down_MMU_BYPASS_TRANSLATION;
      fetch_logic_ctrls_2_up_FetchL1Plugin_logic_WAYS_HIT <= fetch_logic_ctrls_1_down_FetchL1Plugin_logic_WAYS_HIT;
      fetch_logic_ctrls_2_up_GSharePlugin_GSHARE_COUNTER_0 <= fetch_logic_ctrls_1_down_GSharePlugin_GSHARE_COUNTER_0;
      fetch_logic_ctrls_2_up_Prediction_WORD_JUMPED <= fetch_logic_ctrls_1_down_Prediction_WORD_JUMPED;
      fetch_logic_ctrls_2_up_Prediction_WORD_JUMP_PC <= fetch_logic_ctrls_1_down_Prediction_WORD_JUMP_PC;
      fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_BRANCH <= fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_BRANCH;
      fetch_logic_ctrls_2_up_Prediction_WORD_SLICES_TAKEN <= fetch_logic_ctrls_1_down_Prediction_WORD_SLICES_TAKEN;
      fetch_logic_ctrls_2_up_MMU_HAZARD <= fetch_logic_ctrls_1_down_MMU_HAZARD;
      fetch_logic_ctrls_2_up_MMU_REFILL <= fetch_logic_ctrls_1_down_MMU_REFILL;
      fetch_logic_ctrls_2_up_MMU_TRANSLATED <= fetch_logic_ctrls_1_down_MMU_TRANSLATED;
      fetch_logic_ctrls_2_up_MMU_ALLOW_EXECUTE <= fetch_logic_ctrls_1_down_MMU_ALLOW_EXECUTE;
      fetch_logic_ctrls_2_up_MMU_PAGE_FAULT <= fetch_logic_ctrls_1_down_MMU_PAGE_FAULT;
      fetch_logic_ctrls_2_up_MMU_ACCESS_FAULT <= fetch_logic_ctrls_1_down_MMU_ACCESS_FAULT;
    end
    if(decode_ctrls_0_down_isReady) begin
      decode_ctrls_1_up_Decode_INSTRUCTION_0 <= decode_ctrls_0_down_Decode_INSTRUCTION_0;
      decode_ctrls_1_up_Decode_DECOMPRESSION_FAULT_0 <= decode_ctrls_0_down_Decode_DECOMPRESSION_FAULT_0;
      decode_ctrls_1_up_Decode_INSTRUCTION_RAW_0 <= decode_ctrls_0_down_Decode_INSTRUCTION_RAW_0;
      decode_ctrls_1_up_PC_0 <= decode_ctrls_0_down_PC_0;
      decode_ctrls_1_up_Decode_DOP_ID_0 <= decode_ctrls_0_down_Decode_DOP_ID_0;
      decode_ctrls_1_up_GSharePlugin_GSHARE_COUNTER_0_0 <= decode_ctrls_0_down_GSharePlugin_GSHARE_COUNTER_0_0;
      decode_ctrls_1_up_Prediction_BRANCH_HISTORY_0 <= decode_ctrls_0_down_Prediction_BRANCH_HISTORY_0;
      decode_ctrls_1_up_TRAP_0 <= decode_ctrls_0_down_TRAP_0;
      decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_0 <= decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_0;
      decode_ctrls_1_up_Prediction_ALIGNED_JUMPED_PC_0 <= decode_ctrls_0_down_Prediction_ALIGNED_JUMPED_PC_0;
      decode_ctrls_1_up_Prediction_ALIGNED_SLICES_BRANCH_0 <= decode_ctrls_0_down_Prediction_ALIGNED_SLICES_BRANCH_0;
      decode_ctrls_1_up_Prediction_ALIGNED_SLICES_TAKEN_0 <= decode_ctrls_0_down_Prediction_ALIGNED_SLICES_TAKEN_0;
      decode_ctrls_1_up_Prediction_ALIGN_REDO_0 <= decode_ctrls_0_down_Prediction_ALIGN_REDO_0;
    end
    if(execute_ctrl0_down_isReady) begin
      execute_ctrl1_up_Decode_UOP_lane0 <= execute_ctrl0_down_Decode_UOP_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_JUMPED_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_JUMPED_lane0;
      execute_ctrl1_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= execute_ctrl0_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      execute_ctrl1_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= execute_ctrl0_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      execute_ctrl1_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl0_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl1_up_PC_lane0 <= execute_ctrl0_down_PC_lane0;
      execute_ctrl1_up_TRAP_lane0 <= execute_ctrl0_down_TRAP_lane0;
      execute_ctrl1_up_Decode_UOP_ID_lane0 <= execute_ctrl0_down_Decode_UOP_ID_lane0;
      execute_ctrl1_up_RS1_PHYS_lane0 <= execute_ctrl0_down_RS1_PHYS_lane0;
      execute_ctrl1_up_RS2_PHYS_lane0 <= execute_ctrl0_down_RS2_PHYS_lane0;
      execute_ctrl1_up_RD_ENABLE_lane0 <= execute_ctrl0_down_RD_ENABLE_lane0;
      execute_ctrl1_up_RD_PHYS_lane0 <= execute_ctrl0_down_RD_PHYS_lane0;
      execute_ctrl1_up_COMPLETED_lane0 <= execute_ctrl0_down_COMPLETED_lane0;
      execute_ctrl1_up_AguPlugin_SIZE_lane0 <= execute_ctrl0_down_AguPlugin_SIZE_lane0;
    end
    if(execute_ctrl1_down_isReady) begin
      execute_ctrl2_up_Decode_UOP_lane0 <= execute_ctrl1_down_Decode_UOP_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_JUMPED_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_JUMPED_lane0;
      execute_ctrl2_up_Prediction_ALIGNED_JUMPED_PC_lane0 <= execute_ctrl1_down_Prediction_ALIGNED_JUMPED_PC_lane0;
      execute_ctrl2_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= execute_ctrl1_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      execute_ctrl2_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl1_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl2_up_PC_lane0 <= execute_ctrl1_down_PC_lane0;
      execute_ctrl2_up_TRAP_lane0 <= execute_ctrl1_down_TRAP_lane0;
      execute_ctrl2_up_Decode_UOP_ID_lane0 <= execute_ctrl1_down_Decode_UOP_ID_lane0;
      execute_ctrl2_up_RD_ENABLE_lane0 <= execute_ctrl1_down_RD_ENABLE_lane0;
      execute_ctrl2_up_RD_PHYS_lane0 <= execute_ctrl1_down_RD_PHYS_lane0;
      execute_ctrl2_up_COMPLETED_lane0 <= execute_ctrl1_down_COMPLETED_lane0;
      execute_ctrl2_up_AguPlugin_SIZE_lane0 <= execute_ctrl1_down_AguPlugin_SIZE_lane0;
      execute_ctrl2_up_early0_SrcPlugin_SRC1_lane0 <= execute_ctrl1_down_early0_SrcPlugin_SRC1_lane0;
      execute_ctrl2_up_integer_RS1_lane0 <= execute_ctrl1_down_integer_RS1_lane0;
      execute_ctrl2_up_early0_SrcPlugin_SRC2_lane0 <= execute_ctrl1_down_early0_SrcPlugin_SRC2_lane0;
      execute_ctrl2_up_integer_RS2_lane0 <= execute_ctrl1_down_integer_RS2_lane0;
      execute_ctrl2_up_MAY_FLUSH_PRECISE_3_lane0 <= execute_ctrl1_down_MAY_FLUSH_PRECISE_3_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_SEL_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_SEL_lane0;
      execute_ctrl2_up_early0_BarrelShifterPlugin_SEL_lane0 <= execute_ctrl1_down_early0_BarrelShifterPlugin_SEL_lane0;
      execute_ctrl2_up_early0_BranchPlugin_SEL_lane0 <= execute_ctrl1_down_early0_BranchPlugin_SEL_lane0;
      execute_ctrl2_up_early0_MulPlugin_SEL_lane0 <= execute_ctrl1_down_early0_MulPlugin_SEL_lane0;
      execute_ctrl2_up_early0_DivPlugin_SEL_lane0 <= execute_ctrl1_down_early0_DivPlugin_SEL_lane0;
      execute_ctrl2_up_early0_EnvPlugin_SEL_lane0 <= execute_ctrl1_down_early0_EnvPlugin_SEL_lane0;
      execute_ctrl2_up_CfuPlugin_logic_CFU_ENABLE_lane0 <= execute_ctrl1_down_CfuPlugin_logic_CFU_ENABLE_lane0;
      execute_ctrl2_up_CsrAccessPlugin_SEL_lane0 <= execute_ctrl1_down_CsrAccessPlugin_SEL_lane0;
      execute_ctrl2_up_AguPlugin_SEL_lane0 <= execute_ctrl1_down_AguPlugin_SEL_lane0;
      execute_ctrl2_up_LsuPlugin_logic_FENCE_lane0 <= execute_ctrl1_down_LsuPlugin_logic_FENCE_lane0;
      execute_ctrl2_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= execute_ctrl1_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      execute_ctrl2_up_COMPLETION_AT_2_lane0 <= execute_ctrl1_down_COMPLETION_AT_2_lane0;
      execute_ctrl2_up_COMPLETION_AT_3_lane0 <= execute_ctrl1_down_COMPLETION_AT_3_lane0;
      execute_ctrl2_up_COMPLETION_AT_4_lane0 <= execute_ctrl1_down_COMPLETION_AT_4_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_0_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_0_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl2_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl1_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_ALU_ADD_SUB_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_ALU_ADD_SUB_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_ALU_SLTX_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_ALU_SLTX_lane0;
      execute_ctrl2_up_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0 <= execute_ctrl1_down_early0_IntAluPlugin_ALU_BITWISE_CTRL_lane0;
      execute_ctrl2_up_SrcStageables_REVERT_lane0 <= execute_ctrl1_down_SrcStageables_REVERT_lane0;
      execute_ctrl2_up_SrcStageables_ZERO_lane0 <= execute_ctrl1_down_SrcStageables_ZERO_lane0;
      execute_ctrl2_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= execute_ctrl1_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      execute_ctrl2_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= execute_ctrl1_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      execute_ctrl2_up_BYPASSED_AT_3_lane0 <= execute_ctrl1_down_BYPASSED_AT_3_lane0;
      execute_ctrl2_up_SrcStageables_UNSIGNED_lane0 <= execute_ctrl1_down_SrcStageables_UNSIGNED_lane0;
      execute_ctrl2_up_BarrelShifterPlugin_LEFT_lane0 <= execute_ctrl1_down_BarrelShifterPlugin_LEFT_lane0;
      execute_ctrl2_up_BarrelShifterPlugin_SIGNED_lane0 <= execute_ctrl1_down_BarrelShifterPlugin_SIGNED_lane0;
      execute_ctrl2_up_BranchPlugin_BRANCH_CTRL_lane0 <= execute_ctrl1_down_BranchPlugin_BRANCH_CTRL_lane0;
      execute_ctrl2_up_CfuPlugin_logic_CFU_ENCODING_lane0 <= execute_ctrl1_down_CfuPlugin_logic_CFU_ENCODING_lane0;
      execute_ctrl2_up_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0 <= execute_ctrl1_down_CfuPlugin_logic_CFU_INPUT_2_KIND_lane0;
      execute_ctrl2_up_MulPlugin_HIGH_lane0 <= execute_ctrl1_down_MulPlugin_HIGH_lane0;
      execute_ctrl2_up_RsUnsignedPlugin_RS1_SIGNED_lane0 <= execute_ctrl1_down_RsUnsignedPlugin_RS1_SIGNED_lane0;
      execute_ctrl2_up_RsUnsignedPlugin_RS2_SIGNED_lane0 <= execute_ctrl1_down_RsUnsignedPlugin_RS2_SIGNED_lane0;
      execute_ctrl2_up_DivPlugin_REM_lane0 <= execute_ctrl1_down_DivPlugin_REM_lane0;
      execute_ctrl2_up_CsrAccessPlugin_CSR_IMM_lane0 <= execute_ctrl1_down_CsrAccessPlugin_CSR_IMM_lane0;
      execute_ctrl2_up_CsrAccessPlugin_CSR_MASK_lane0 <= execute_ctrl1_down_CsrAccessPlugin_CSR_MASK_lane0;
      execute_ctrl2_up_CsrAccessPlugin_CSR_CLEAR_lane0 <= execute_ctrl1_down_CsrAccessPlugin_CSR_CLEAR_lane0;
      execute_ctrl2_up_AguPlugin_LOAD_lane0 <= execute_ctrl1_down_AguPlugin_LOAD_lane0;
      execute_ctrl2_up_AguPlugin_STORE_lane0 <= execute_ctrl1_down_AguPlugin_STORE_lane0;
      execute_ctrl2_up_AguPlugin_ATOMIC_lane0 <= execute_ctrl1_down_AguPlugin_ATOMIC_lane0;
      execute_ctrl2_up_AguPlugin_FLOAT_lane0 <= execute_ctrl1_down_AguPlugin_FLOAT_lane0;
      execute_ctrl2_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= execute_ctrl1_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      execute_ctrl2_up_early0_EnvPlugin_OP_lane0 <= execute_ctrl1_down_early0_EnvPlugin_OP_lane0;
    end
    if(execute_ctrl2_down_isReady) begin
      execute_ctrl3_up_Decode_UOP_lane0 <= execute_ctrl2_down_Decode_UOP_lane0;
      execute_ctrl3_up_Prediction_ALIGNED_JUMPED_lane0 <= execute_ctrl2_down_Prediction_ALIGNED_JUMPED_lane0;
      execute_ctrl3_up_GSharePlugin_GSHARE_COUNTER_lane0_0 <= execute_ctrl2_down_GSharePlugin_GSHARE_COUNTER_lane0_0;
      execute_ctrl3_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl2_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl3_up_PC_lane0 <= execute_ctrl2_down_PC_lane0;
      execute_ctrl3_up_TRAP_lane0 <= execute_ctrl2_down_TRAP_lane0;
      execute_ctrl3_up_Decode_UOP_ID_lane0 <= execute_ctrl2_down_Decode_UOP_ID_lane0;
      execute_ctrl3_up_RD_ENABLE_lane0 <= execute_ctrl2_down_RD_ENABLE_lane0;
      execute_ctrl3_up_RD_PHYS_lane0 <= execute_ctrl2_down_RD_PHYS_lane0;
      execute_ctrl3_up_COMPLETED_lane0 <= execute_ctrl2_down_COMPLETED_lane0;
      execute_ctrl3_up_AguPlugin_SIZE_lane0 <= execute_ctrl2_down_AguPlugin_SIZE_lane0;
      execute_ctrl3_up_integer_RS2_lane0 <= execute_ctrl2_down_integer_RS2_lane0;
      execute_ctrl3_up_early0_BranchPlugin_SEL_lane0 <= execute_ctrl2_down_early0_BranchPlugin_SEL_lane0;
      execute_ctrl3_up_early0_MulPlugin_SEL_lane0 <= execute_ctrl2_down_early0_MulPlugin_SEL_lane0;
      execute_ctrl3_up_early0_DivPlugin_SEL_lane0 <= execute_ctrl2_down_early0_DivPlugin_SEL_lane0;
      execute_ctrl3_up_CfuPlugin_logic_CFU_ENABLE_lane0 <= execute_ctrl2_down_CfuPlugin_logic_CFU_ENABLE_lane0;
      execute_ctrl3_up_CsrAccessPlugin_SEL_lane0 <= execute_ctrl2_down_CsrAccessPlugin_SEL_lane0;
      execute_ctrl3_up_AguPlugin_SEL_lane0 <= execute_ctrl2_down_AguPlugin_SEL_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FENCE_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FENCE_lane0;
      execute_ctrl3_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= execute_ctrl2_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      execute_ctrl3_up_COMPLETION_AT_3_lane0 <= execute_ctrl2_down_COMPLETION_AT_3_lane0;
      execute_ctrl3_up_COMPLETION_AT_4_lane0 <= execute_ctrl2_down_COMPLETION_AT_4_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_1_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_1_ENABLE_lane0;
      execute_ctrl3_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl2_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl3_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= execute_ctrl2_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      execute_ctrl3_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= execute_ctrl2_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      execute_ctrl3_up_BranchPlugin_BRANCH_CTRL_lane0 <= execute_ctrl2_down_BranchPlugin_BRANCH_CTRL_lane0;
      execute_ctrl3_up_MulPlugin_HIGH_lane0 <= execute_ctrl2_down_MulPlugin_HIGH_lane0;
      execute_ctrl3_up_AguPlugin_LOAD_lane0 <= execute_ctrl2_down_AguPlugin_LOAD_lane0;
      execute_ctrl3_up_AguPlugin_STORE_lane0 <= execute_ctrl2_down_AguPlugin_STORE_lane0;
      execute_ctrl3_up_AguPlugin_ATOMIC_lane0 <= execute_ctrl2_down_AguPlugin_ATOMIC_lane0;
      execute_ctrl3_up_AguPlugin_FLOAT_lane0 <= execute_ctrl2_down_AguPlugin_FLOAT_lane0;
      execute_ctrl3_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= execute_ctrl2_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      execute_ctrl3_up_COMMIT_lane0 <= execute_ctrl2_down_COMMIT_lane0;
      execute_ctrl3_up_early0_SrcPlugin_ADD_SUB_lane0 <= execute_ctrl2_down_early0_SrcPlugin_ADD_SUB_lane0;
      execute_ctrl3_up_early0_SrcPlugin_LESS_lane0 <= execute_ctrl2_down_early0_SrcPlugin_LESS_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_0_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_1_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_2_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
      execute_ctrl3_up_early0_MulPlugin_logic_mul_VALUES_3_lane0 <= execute_ctrl2_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
      execute_ctrl3_up_DivPlugin_DIV_RESULT_lane0 <= execute_ctrl2_down_DivPlugin_DIV_RESULT_lane0;
      execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_TRUE_lane0 <= execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_TRUE_lane0;
      execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_FALSE_lane0 <= execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_FALSE_lane0;
      execute_ctrl3_up_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0 <= execute_ctrl2_down_early0_BranchPlugin_pcCalc_PC_LAST_SLICE_lane0;
      execute_ctrl3_up_early0_BranchPlugin_logic_alu_EQ_lane0 <= execute_ctrl2_down_early0_BranchPlugin_logic_alu_EQ_lane0;
      execute_ctrl3_up_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0 <= execute_ctrl2_down_early0_BranchPlugin_logic_alu_btb_BAD_TARGET_lane0;
      execute_ctrl3_up_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0 <= execute_ctrl2_down_early0_BranchPlugin_logic_alu_MSB_FAILED_lane0;
      execute_ctrl3_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl2_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      execute_ctrl3_up_LsuL1_MIXED_ADDRESS_lane0 <= execute_ctrl2_down_LsuL1_MIXED_ADDRESS_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_BANK_BUSY_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_BANK_BUSY_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_VALID_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_ADDRESS_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALID_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0 <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_0;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_1 <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_plru_1;
      execute_ctrl3_up_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty <= execute_ctrl2_down_LsuL1Plugin_logic_lsu_rt0_SHARED_BYPASS_VALUE_lane0_dirty;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
      execute_ctrl3_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 <= execute_ctrl2_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FORCE_PHYSICAL_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FORCE_PHYSICAL_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_ACCESS_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_ACCESS_lane0;
      execute_ctrl3_up_LsuL1_MASK_lane0 <= execute_ctrl2_down_LsuL1_MASK_lane0;
      execute_ctrl3_up_LsuL1_SIZE_lane0 <= execute_ctrl2_down_LsuL1_SIZE_lane0;
      execute_ctrl3_up_LsuL1_LOAD_lane0 <= execute_ctrl2_down_LsuL1_LOAD_lane0;
      execute_ctrl3_up_LsuL1_ATOMIC_lane0 <= execute_ctrl2_down_LsuL1_ATOMIC_lane0;
      execute_ctrl3_up_LsuL1_STORE_lane0 <= execute_ctrl2_down_LsuL1_STORE_lane0;
      execute_ctrl3_up_LsuL1_CLEAN_lane0 <= execute_ctrl2_down_LsuL1_CLEAN_lane0;
      execute_ctrl3_up_LsuL1_INVALID_lane0 <= execute_ctrl2_down_LsuL1_INVALID_lane0;
      execute_ctrl3_up_LsuL1_PREFETCH_lane0 <= execute_ctrl2_down_LsuL1_PREFETCH_lane0;
      execute_ctrl3_up_LsuL1_FLUSH_lane0 <= execute_ctrl2_down_LsuL1_FLUSH_lane0;
      execute_ctrl3_up_Decode_STORE_ID_lane0 <= execute_ctrl2_down_Decode_STORE_ID_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_LSU_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_LSU_lane0;
      execute_ctrl3_up_LsuPlugin_logic_FROM_PREFETCH_lane0 <= execute_ctrl2_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_valid <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_valid;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_virtualAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_virtualAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_physicalAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_physicalAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowRead <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowRead;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowWrite <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowWrite;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowExecute <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowExecute;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_0_allowUser <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_0_allowUser;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_valid <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_valid;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_virtualAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_virtualAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_physicalAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_physicalAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowRead <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowRead;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowWrite <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowWrite;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowExecute <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowExecute;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_1_allowUser <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_1_allowUser;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_valid <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_valid;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_virtualAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_virtualAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_physicalAddress <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_physicalAddress;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowRead <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowRead;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowWrite <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowWrite;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowExecute <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowExecute;
      execute_ctrl3_up_MMU_L0_ENTRIES_lane0_2_allowUser <= execute_ctrl2_down_MMU_L0_ENTRIES_lane0_2_allowUser;
      execute_ctrl3_up_MMU_L0_HITS_PRE_VALID_lane0 <= execute_ctrl2_down_MMU_L0_HITS_PRE_VALID_lane0;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_valid <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_valid;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_virtualAddress <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_virtualAddress;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_physicalAddress <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_physicalAddress;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowRead <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowRead;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowWrite <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowWrite;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowExecute <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowExecute;
      execute_ctrl3_up_MMU_L1_ENTRIES_lane0_0_allowUser <= execute_ctrl2_down_MMU_L1_ENTRIES_lane0_0_allowUser;
      execute_ctrl3_up_MMU_L1_HITS_PRE_VALID_lane0 <= execute_ctrl2_down_MMU_L1_HITS_PRE_VALID_lane0;
    end
    if(execute_ctrl3_down_isReady) begin
      execute_ctrl4_up_Decode_UOP_lane0 <= execute_ctrl3_down_Decode_UOP_lane0;
      execute_ctrl4_up_Prediction_BRANCH_HISTORY_lane0 <= execute_ctrl3_down_Prediction_BRANCH_HISTORY_lane0;
      execute_ctrl4_up_PC_lane0 <= execute_ctrl3_down_PC_lane0;
      execute_ctrl4_up_TRAP_lane0 <= execute_ctrl3_down_TRAP_lane0;
      execute_ctrl4_up_Decode_UOP_ID_lane0 <= execute_ctrl3_down_Decode_UOP_ID_lane0;
      execute_ctrl4_up_RD_ENABLE_lane0 <= execute_ctrl3_down_RD_ENABLE_lane0;
      execute_ctrl4_up_RD_PHYS_lane0 <= execute_ctrl3_down_RD_PHYS_lane0;
      execute_ctrl4_up_COMPLETED_lane0 <= execute_ctrl3_down_COMPLETED_lane0;
      execute_ctrl4_up_AguPlugin_SIZE_lane0 <= execute_ctrl3_down_AguPlugin_SIZE_lane0;
      execute_ctrl4_up_integer_RS2_lane0 <= execute_ctrl3_down_integer_RS2_lane0;
      execute_ctrl4_up_early0_MulPlugin_SEL_lane0 <= execute_ctrl3_down_early0_MulPlugin_SEL_lane0;
      execute_ctrl4_up_CfuPlugin_logic_CFU_ENABLE_lane0 <= execute_ctrl3_down_CfuPlugin_logic_CFU_ENABLE_lane0;
      execute_ctrl4_up_AguPlugin_SEL_lane0 <= execute_ctrl3_down_AguPlugin_SEL_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FENCE_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FENCE_lane0;
      execute_ctrl4_up_lane0_integer_WriteBackPlugin_SEL_lane0 <= execute_ctrl3_down_lane0_integer_WriteBackPlugin_SEL_lane0;
      execute_ctrl4_up_COMPLETION_AT_4_lane0 <= execute_ctrl3_down_COMPLETION_AT_4_lane0;
      execute_ctrl4_up_lane0_logic_completions_onCtrl_2_ENABLE_lane0 <= execute_ctrl3_down_lane0_logic_completions_onCtrl_2_ENABLE_lane0;
      execute_ctrl4_up_lane0_IntFormatPlugin_logic_SIGNED_lane0 <= execute_ctrl3_down_lane0_IntFormatPlugin_logic_SIGNED_lane0;
      execute_ctrl4_up_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0 <= execute_ctrl3_down_lane0_IntFormatPlugin_logic_WIDTH_ID_lane0;
      execute_ctrl4_up_MulPlugin_HIGH_lane0 <= execute_ctrl3_down_MulPlugin_HIGH_lane0;
      execute_ctrl4_up_AguPlugin_LOAD_lane0 <= execute_ctrl3_down_AguPlugin_LOAD_lane0;
      execute_ctrl4_up_AguPlugin_STORE_lane0 <= execute_ctrl3_down_AguPlugin_STORE_lane0;
      execute_ctrl4_up_AguPlugin_ATOMIC_lane0 <= execute_ctrl3_down_AguPlugin_ATOMIC_lane0;
      execute_ctrl4_up_AguPlugin_FLOAT_lane0 <= execute_ctrl3_down_AguPlugin_FLOAT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_LSU_PREFETCH_lane0 <= execute_ctrl3_down_LsuPlugin_logic_LSU_PREFETCH_lane0;
      execute_ctrl4_up_COMMIT_lane0 <= execute_ctrl3_down_COMMIT_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_0_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_0_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_1_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_1_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_2_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_2_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_mul_VALUES_3_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_mul_VALUES_3_lane0;
      execute_ctrl4_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl3_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
      execute_ctrl4_up_LsuL1_MIXED_ADDRESS_lane0 <= execute_ctrl3_down_LsuL1_MIXED_ADDRESS_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_DATA_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_EVENT_WRITE_MASK_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FROM_ACCESS_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FROM_ACCESS_lane0;
      execute_ctrl4_up_LsuL1_MASK_lane0 <= execute_ctrl3_down_LsuL1_MASK_lane0;
      execute_ctrl4_up_LsuL1_SIZE_lane0 <= execute_ctrl3_down_LsuL1_SIZE_lane0;
      execute_ctrl4_up_LsuL1_LOAD_lane0 <= execute_ctrl3_down_LsuL1_LOAD_lane0;
      execute_ctrl4_up_LsuL1_ATOMIC_lane0 <= execute_ctrl3_down_LsuL1_ATOMIC_lane0;
      execute_ctrl4_up_LsuL1_STORE_lane0 <= execute_ctrl3_down_LsuL1_STORE_lane0;
      execute_ctrl4_up_LsuL1_CLEAN_lane0 <= execute_ctrl3_down_LsuL1_CLEAN_lane0;
      execute_ctrl4_up_LsuL1_INVALID_lane0 <= execute_ctrl3_down_LsuL1_INVALID_lane0;
      execute_ctrl4_up_LsuL1_PREFETCH_lane0 <= execute_ctrl3_down_LsuL1_PREFETCH_lane0;
      execute_ctrl4_up_LsuL1_FLUSH_lane0 <= execute_ctrl3_down_LsuL1_FLUSH_lane0;
      execute_ctrl4_up_Decode_STORE_ID_lane0 <= execute_ctrl3_down_Decode_STORE_ID_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FROM_LSU_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FROM_LSU_lane0;
      execute_ctrl4_up_LsuPlugin_logic_FROM_PREFETCH_lane0 <= execute_ctrl3_down_LsuPlugin_logic_FROM_PREFETCH_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_0 <= execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_0;
      execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_plru_1 <= execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_plru_1;
      execute_ctrl4_up_LsuL1Plugin_logic_SHARED_lane0_dirty <= execute_ctrl3_down_LsuL1Plugin_logic_SHARED_lane0_dirty;
      execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_0_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_0_lane0;
      execute_ctrl4_up_early0_MulPlugin_logic_steps_0_adders_1_lane0 <= execute_ctrl3_down_early0_MulPlugin_logic_steps_0_adders_1_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_BANK_BUSY_REMAPPED_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_0 <= execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_0;
      execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_1 <= execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_1;
      execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_2 <= execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_2;
      execute_ctrl4_up_LsuL1Plugin_logic_BANKS_MUXES_lane0_3 <= execute_ctrl3_down_LsuL1Plugin_logic_BANKS_MUXES_lane0_3;
      execute_ctrl4_up_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_WRITE_TO_READ_HAZARDS_lane0;
      execute_ctrl4_up_LsuL1_PHYSICAL_ADDRESS_lane0 <= execute_ctrl3_down_LsuL1_PHYSICAL_ADDRESS_lane0;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_loaded;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_address;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_0_fault;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_loaded;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_address;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_1_fault;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_loaded;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_address;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_2_fault;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_loaded;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_address;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_TAGS_lane0_3_fault;
      execute_ctrl4_up_LsuL1Plugin_logic_WAYS_HITS_lane0 <= execute_ctrl3_down_LsuL1Plugin_logic_WAYS_HITS_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onTrigger_HIT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onTrigger_HIT_lane0;
      execute_ctrl4_up_MMU_TRANSLATED_lane0 <= execute_ctrl3_down_MMU_TRANSLATED_lane0;
      execute_ctrl4_up_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0 <= execute_ctrl3_down_LsuPlugin_logic_preCtrl_MISS_ALIGNED_lane0;
      execute_ctrl4_up_LsuPlugin_logic_preCtrl_IS_AMO_lane0 <= execute_ctrl3_down_LsuPlugin_logic_preCtrl_IS_AMO_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault <= execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_fault;
      execute_ctrl4_up_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io <= execute_ctrl3_down_LsuPlugin_logic_onPma_CACHED_RSP_lane0_io;
      execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_fault <= execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_fault;
      execute_ctrl4_up_LsuPlugin_logic_onPma_IO_RSP_lane0_io <= execute_ctrl3_down_LsuPlugin_logic_onPma_IO_RSP_lane0_io;
      execute_ctrl4_up_LsuPlugin_logic_onPma_IO_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onPma_IO_lane0;
      execute_ctrl4_up_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0 <= execute_ctrl3_down_LsuPlugin_logic_onPma_FROM_LSU_MSB_FAILED_lane0;
      execute_ctrl4_up_LsuPlugin_logic_MMU_PAGE_FAULT_lane0 <= execute_ctrl3_down_LsuPlugin_logic_MMU_PAGE_FAULT_lane0;
      execute_ctrl4_up_LsuPlugin_logic_MMU_FAILURE_lane0 <= execute_ctrl3_down_LsuPlugin_logic_MMU_FAILURE_lane0;
      execute_ctrl4_up_MMU_ACCESS_FAULT_lane0 <= execute_ctrl3_down_MMU_ACCESS_FAULT_lane0;
      execute_ctrl4_up_MMU_REFILL_lane0 <= execute_ctrl3_down_MMU_REFILL_lane0;
      execute_ctrl4_up_MMU_HAZARD_lane0 <= execute_ctrl3_down_MMU_HAZARD_lane0;
      execute_ctrl4_up_MMU_BYPASS_TRANSLATION_lane0 <= execute_ctrl3_down_MMU_BYPASS_TRANSLATION_lane0;
    end
    if(execute_ctrl4_down_isReady) begin
      execute_ctrl5_up_RD_ENABLE_lane0 <= execute_ctrl4_down_RD_ENABLE_lane0;
      execute_ctrl5_up_RD_PHYS_lane0 <= execute_ctrl4_down_RD_PHYS_lane0;
      execute_ctrl5_up_COMMIT_lane0 <= execute_ctrl4_down_COMMIT_lane0;
      execute_ctrl5_up_lane0_integer_WriteBackPlugin_logic_DATA_lane0 <= execute_ctrl4_down_lane0_integer_WriteBackPlugin_logic_DATA_lane0;
    end
    case(LsuPlugin_logic_flusher_stateReg)
      LsuPlugin_logic_flusher_CMD : begin
        if(when_LsuPlugin_l363) begin
          LsuPlugin_logic_flusher_waiter <= LsuL1_WRITEBACK_BUSY;
        end
      end
      LsuPlugin_logic_flusher_COMPLETION : begin
        LsuPlugin_logic_flusher_waiter <= (LsuPlugin_logic_flusher_waiter & LsuL1_WRITEBACK_BUSY);
      end
      default : begin
        LsuPlugin_logic_flusher_cmdCounter <= 7'h0;
      end
    endcase
    case(TrapPlugin_logic_harts_0_trap_fsm_stateReg)
      TrapPlugin_logic_harts_0_trap_fsm_RUNNING : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_PROCESS_1 : begin
        TrapPlugin_logic_harts_0_trap_fsm_triggerEbreakReg <= TrapPlugin_logic_harts_0_trap_fsm_triggerEbreak;
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVAL : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_TVEC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_TRAP_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_EPC : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_XRET_APPLY : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_ATS_RSP : begin
        if(TrapPlugin_logic_harts_0_trap_fsm_atsPorts_refill_rsp_valid) begin
          if(when_TrapPlugin_l509) begin
            TrapPlugin_logic_harts_0_trap_pending_state_exception <= 1'b1;
            case(switch_TrapPlugin_l511)
              3'b110 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b0001;
              end
              3'b100 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b0101;
              end
              3'b101 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b0111;
              end
              3'b010 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b1100;
              end
              3'b000 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b1101;
              end
              3'b001 : begin
                TrapPlugin_logic_harts_0_trap_pending_state_code <= 4'b1111;
              end
              default : begin
              end
            endcase
          end
        end
      end
      TrapPlugin_logic_harts_0_trap_fsm_JUMP : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_LSU_FLUSH : begin
      end
      TrapPlugin_logic_harts_0_trap_fsm_FETCH_FLUSH : begin
      end
      default : begin
      end
    endcase
    case(MmuPlugin_logic_refill_stateReg)
      MmuPlugin_logic_refill_IDLE : begin
        if(MmuPlugin_logic_refill_arbiter_io_output_valid) begin
          MmuPlugin_logic_refill_portOhReg <= MmuPlugin_logic_refill_arbiter_io_chosenOH;
          MmuPlugin_logic_refill_storageOhReg <= (2'b01 <<< MmuPlugin_logic_refill_arbiter_io_output_payload_storageId);
          MmuPlugin_logic_refill_virtual <= MmuPlugin_logic_refill_arbiter_io_output_payload_address;
          MmuPlugin_logic_refill_load_address <= {{MmuPlugin_logic_satp_ppn,MmuPlugin_logic_refill_arbiter_io_output_payload_address[31 : 22]},2'b00};
        end
      end
      MmuPlugin_logic_refill_CMD_0 : begin
      end
      MmuPlugin_logic_refill_CMD_1 : begin
      end
      MmuPlugin_logic_refill_RSP_0 : begin
      end
      MmuPlugin_logic_refill_RSP_1 : begin
        if(MmuPlugin_logic_refill_load_rsp_valid) begin
          if(!MmuPlugin_logic_refill_load_rsp_payload_redo) begin
            if(!when_MmuPlugin_l487) begin
              MmuPlugin_logic_refill_load_address <= MmuPlugin_logic_refill_load_nextLevelBase;
              MmuPlugin_logic_refill_load_address[11 : 2] <= MmuPlugin_logic_refill_virtual[21 : 12];
            end
          end
        end
      end
      default : begin
      end
    endcase
    case(PerformanceCounterPlugin_logic_fsm_stateReg)
      PerformanceCounterPlugin_logic_fsm_IDLE : begin
        PerformanceCounterPlugin_logic_fsm_cmd_oh <= {(PerformanceCounterPlugin_logic_fsm_idleCsrAddress == 2'b10),(PerformanceCounterPlugin_logic_fsm_idleCsrAddress == 2'b00)};
        if(!PerformanceCounterPlugin_logic_fsm_csrWriteCmd_valid) begin
          if(PerformanceCounterPlugin_logic_fsm_flusherCmd_valid) begin
            PerformanceCounterPlugin_logic_fsm_cmd_flusher <= 1'b1;
            PerformanceCounterPlugin_logic_fsm_cmd_oh <= PerformanceCounterPlugin_logic_fsm_flusherCmd_payload_oh;
          end else begin
            if(PerformanceCounterPlugin_logic_fsm_csrReadCmd_valid) begin
              PerformanceCounterPlugin_logic_fsm_cmd_flusher <= 1'b0;
            end
          end
        end
        PerformanceCounterPlugin_logic_fsm_carry <= 1'b0;
      end
      PerformanceCounterPlugin_logic_fsm_READ_LOW : begin
        PerformanceCounterPlugin_logic_fsm_ramReaded <= PerformanceCounterPlugin_logic_readPort_data;
        PerformanceCounterPlugin_logic_fsm_counterReaded <= ((_zz_PerformanceCounterPlugin_logic_fsm_cmd_address ? PerformanceCounterPlugin_logic_counters_cycle_value : 8'h0) | (_zz_PerformanceCounterPlugin_logic_fsm_cmd_address_1 ? PerformanceCounterPlugin_logic_counters_instret_value : 8'h0));
      end
      PerformanceCounterPlugin_logic_fsm_CALC_LOW : begin
        if(PerformanceCounterPlugin_logic_writePort_ready) begin
          if(when_PerformanceCounterPlugin_l278) begin
            PerformanceCounterPlugin_logic_fsm_carry <= 1'b1;
          end
        end
      end
      PerformanceCounterPlugin_logic_fsm_READ_HIGH : begin
        PerformanceCounterPlugin_logic_fsm_ramReaded <= PerformanceCounterPlugin_logic_readPort_data;
      end
      PerformanceCounterPlugin_logic_fsm_CALC_HIGH : begin
      end
      PerformanceCounterPlugin_logic_fsm_CSR_WRITE : begin
      end
      default : begin
      end
    endcase
    case(CsrAccessPlugin_logic_fsm_stateReg)
      CsrAccessPlugin_logic_fsm_READ : begin
        CsrAccessPlugin_logic_fsm_interface_aluInput <= CsrAccessPlugin_bus_read_toWriteBits;
        CsrAccessPlugin_logic_fsm_interface_csrValue <= CsrAccessPlugin_logic_fsm_readLogic_csrValue;
      end
      CsrAccessPlugin_logic_fsm_WRITE : begin
      end
      CsrAccessPlugin_logic_fsm_COMPLETION : begin
      end
      default : begin
        REG_CSR_768 <= COMB_CSR_768;
        REG_CSR_256 <= COMB_CSR_256;
        REG_CSR_384 <= COMB_CSR_384;
        REG_CSR_3008 <= COMB_CSR_3008;
        REG_CSR_1952 <= COMB_CSR_1952;
        REG_CSR_1953 <= COMB_CSR_1953;
        REG_CSR_1954 <= COMB_CSR_1954;
        REG_CSR_3857 <= COMB_CSR_3857;
        REG_CSR_3858 <= COMB_CSR_3858;
        REG_CSR_3859 <= COMB_CSR_3859;
        REG_CSR_3860 <= COMB_CSR_3860;
        REG_CSR_769 <= COMB_CSR_769;
        REG_CSR_834 <= COMB_CSR_834;
        REG_CSR_836 <= COMB_CSR_836;
        REG_CSR_772 <= COMB_CSR_772;
        REG_CSR_770 <= COMB_CSR_770;
        REG_CSR_771 <= COMB_CSR_771;
        REG_CSR_322 <= COMB_CSR_322;
        REG_CSR_260 <= COMB_CSR_260;
        REG_CSR_324 <= COMB_CSR_324;
        REG_CSR_3073 <= COMB_CSR_3073;
        REG_CSR_3201 <= COMB_CSR_3201;
        REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter <= COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_tvecFilter;
        REG_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter <= COMB_CSR_PrivilegedPlugin_logic_readAnyWriteLegal_epcFilter;
        REG_CSR_774 <= COMB_CSR_774;
        REG_CSR_262 <= COMB_CSR_262;
        REG_CSR_800 <= COMB_CSR_800;
        REG_CSR_ <= COMB_CSR_;
        REG_CSR_CsrRamPlugin_csrMapper_selFilter <= COMB_CSR_CsrRamPlugin_csrMapper_selFilter;
        REG_CSR_PerformanceCounterPlugin_logic_csrFilter <= COMB_CSR_PerformanceCounterPlugin_logic_csrFilter;
        REG_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter <= COMB_CSR_CsrAccessPlugin_logic_trapNextOnWriteFilter;
      end
    endcase
  end


endmodule

module StreamArbiter_9 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_opcode,
  input  wire [2:0]    io_inputs_0_payload_param,
  input  wire [2:0]    io_inputs_0_payload_source,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire          io_inputs_0_payload_denied,
  input  wire [31:0]   io_inputs_0_payload_data,
  input  wire          io_inputs_0_payload_corrupt,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_opcode,
  input  wire [2:0]    io_inputs_1_payload_param,
  input  wire [2:0]    io_inputs_1_payload_source,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire          io_inputs_1_payload_denied,
  input  wire [31:0]   io_inputs_1_payload_data,
  input  wire          io_inputs_1_payload_corrupt,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [2:0]    io_inputs_2_payload_opcode,
  input  wire [2:0]    io_inputs_2_payload_param,
  input  wire [2:0]    io_inputs_2_payload_source,
  input  wire [2:0]    io_inputs_2_payload_size,
  input  wire          io_inputs_2_payload_denied,
  input  wire [31:0]   io_inputs_2_payload_data,
  input  wire          io_inputs_2_payload_corrupt,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_opcode,
  output wire [2:0]    io_output_payload_param,
  output wire [2:0]    io_output_payload_source,
  output wire [2:0]    io_output_payload_size,
  output wire          io_output_payload_denied,
  output wire [31:0]   io_output_payload_data,
  output wire          io_output_payload_corrupt,
  output wire [1:0]    io_chosen,
  output wire [2:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          litex_reset
);
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire       [5:0]    _zz__zz_maskProposal_0_2;
  wire       [5:0]    _zz__zz_maskProposal_0_2_1;
  wire       [2:0]    _zz__zz_maskProposal_0_2_2;
  reg        [3:0]    _zz_io_output_tracker_last;
  reg        [2:0]    _zz__zz_io_output_payload_opcode;
  reg        [2:0]    _zz_io_output_payload_param_1;
  reg        [2:0]    _zz_io_output_payload_source;
  reg        [2:0]    _zz_io_output_payload_size;
  reg                 _zz_io_output_payload_denied;
  reg        [31:0]   _zz_io_output_payload_data;
  reg                 _zz_io_output_payload_corrupt;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire       [2:0]    _zz_maskProposal_0;
  wire       [5:0]    _zz_maskProposal_0_1;
  wire       [5:0]    _zz_maskProposal_0_2;
  wire       [2:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  reg        [3:0]    io_output_tracker_beat;
  wire                io_output_tracker_last;
  wire                when_Stream_l800;
  wire       [1:0]    _zz_io_output_payload_param;
  wire       [2:0]    _zz_io_output_payload_opcode;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  `ifndef SYNTHESIS
  reg [119:0] io_inputs_0_payload_opcode_string;
  reg [119:0] io_inputs_1_payload_opcode_string;
  reg [119:0] io_inputs_2_payload_opcode_string;
  reg [119:0] io_output_payload_opcode_string;
  reg [119:0] _zz_io_output_payload_opcode_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_1,{maskLocked_0,maskLocked_2}};
  assign _zz__zz_maskProposal_0_2_1 = {3'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(io_output_payload_size)
      3'b000 : _zz_io_output_tracker_last = 4'b0000;
      3'b001 : _zz_io_output_tracker_last = 4'b0000;
      3'b010 : _zz_io_output_tracker_last = 4'b0000;
      3'b011 : _zz_io_output_tracker_last = 4'b0001;
      3'b100 : _zz_io_output_tracker_last = 4'b0011;
      3'b101 : _zz_io_output_tracker_last = 4'b0111;
      default : _zz_io_output_tracker_last = 4'b1111;
    endcase
  end

  always @(*) begin
    case(_zz_io_output_payload_param)
      2'b00 : begin
        _zz__zz_io_output_payload_opcode = io_inputs_0_payload_opcode;
        _zz_io_output_payload_param_1 = io_inputs_0_payload_param;
        _zz_io_output_payload_source = io_inputs_0_payload_source;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_denied = io_inputs_0_payload_denied;
        _zz_io_output_payload_data = io_inputs_0_payload_data;
        _zz_io_output_payload_corrupt = io_inputs_0_payload_corrupt;
      end
      2'b01 : begin
        _zz__zz_io_output_payload_opcode = io_inputs_1_payload_opcode;
        _zz_io_output_payload_param_1 = io_inputs_1_payload_param;
        _zz_io_output_payload_source = io_inputs_1_payload_source;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_denied = io_inputs_1_payload_denied;
        _zz_io_output_payload_data = io_inputs_1_payload_data;
        _zz_io_output_payload_corrupt = io_inputs_1_payload_corrupt;
      end
      default : begin
        _zz__zz_io_output_payload_opcode = io_inputs_2_payload_opcode;
        _zz_io_output_payload_param_1 = io_inputs_2_payload_param;
        _zz_io_output_payload_source = io_inputs_2_payload_source;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_denied = io_inputs_2_payload_denied;
        _zz_io_output_payload_data = io_inputs_2_payload_data;
        _zz_io_output_payload_corrupt = io_inputs_2_payload_corrupt;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_opcode)
      D_ACCESS_ACK : io_inputs_0_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_inputs_0_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_inputs_0_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_inputs_0_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_inputs_0_payload_opcode_string = "RELEASE_ACK    ";
      default : io_inputs_0_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_opcode)
      D_ACCESS_ACK : io_inputs_1_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_inputs_1_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_inputs_1_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_inputs_1_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_inputs_1_payload_opcode_string = "RELEASE_ACK    ";
      default : io_inputs_1_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_opcode)
      D_ACCESS_ACK : io_inputs_2_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_inputs_2_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_inputs_2_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_inputs_2_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_inputs_2_payload_opcode_string = "RELEASE_ACK    ";
      default : io_inputs_2_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_opcode)
      D_ACCESS_ACK : io_output_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_output_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_output_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_output_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_output_payload_opcode_string = "RELEASE_ACK    ";
      default : io_output_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_opcode)
      D_ACCESS_ACK : _zz_io_output_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_output_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_output_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_output_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_output_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_output_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign _zz_maskProposal_0 = {io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[5 : 3] | _zz_maskProposal_0_2[2 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign maskProposal_2 = _zz_maskProposal_0_3[2];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_tracker_last = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_output_payload_opcode)) || (D_GRANT_DATA == io_output_payload_opcode))) || (io_output_tracker_beat == _zz_io_output_tracker_last));
  assign when_Stream_l800 = (io_output_fire && io_output_tracker_last);
  assign io_output_valid = (((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2));
  assign _zz_io_output_payload_param = {maskRouted_2,maskRouted_1};
  assign _zz_io_output_payload_opcode = _zz__zz_io_output_payload_opcode;
  assign io_output_payload_opcode = _zz_io_output_payload_opcode;
  assign io_output_payload_param = _zz_io_output_payload_param_1;
  assign io_output_payload_source = _zz_io_output_payload_source;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_denied = _zz_io_output_payload_denied;
  assign io_output_payload_data = _zz_io_output_payload_data;
  assign io_output_payload_corrupt = _zz_io_output_payload_corrupt;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_chosenOH = {maskRouted_2,{maskRouted_1,maskRouted_0}};
  assign _zz_io_chosen = io_chosenOH[1];
  assign _zz_io_chosen_1 = io_chosenOH[2];
  assign io_chosen = {_zz_io_chosen_1,_zz_io_chosen};
  always @(posedge litex_clk or posedge litex_reset) begin
    if(litex_reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b0;
      maskLocked_2 <= 1'b1;
      io_output_tracker_beat <= 4'b0000;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
        maskLocked_2 <= maskRouted_2;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        io_output_tracker_beat <= (io_output_tracker_beat + 4'b0001);
        if(io_output_tracker_last) begin
          io_output_tracker_beat <= 4'b0000;
        end
      end
      if(when_Stream_l800) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module ContextAsyncBufferFull_1 (
  input  wire          io_add_valid,
  output wire          io_add_ready,
  input  wire [1:0]    io_add_payload_id,
  input  wire [0:0]    io_add_payload_context,
  input  wire          io_remove_valid,
  input  wire [1:0]    io_remove_payload_id,
  input  wire [1:0]    io_query_id,
  output wire [0:0]    io_query_context,
  input  wire          litex_clk
);

  wire                contexts_wr_en;
  wire       [0:0]    contexts_wr_data;
  wire       [0:0]    contexts_rd_data;
  reg                 _zz_wr_en;
  wire                write_valid;
  wire       [1:0]    write_payload_address;
  wire       [0:0]    write_payload_data;
  wire       [1:0]    read_address;
  wire       [0:0]    read_data;

  Ram_1w_1ra #(
    .wordCount      (4         ),
    .wordWidth      (1         ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (2         ),
    .wrDataWidth    (1         ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (2         ),
    .rdDataWidth    (1         )
  ) contexts (
    .clk     (litex_clk                 ), //i
    .wr_en   (contexts_wr_en            ), //i
    .wr_mask (1'b1                      ), //i
    .wr_addr (write_payload_address[1:0]), //i
    .wr_data (contexts_wr_data          ), //i
    .rd_addr (read_address[1:0]         ), //i
    .rd_data (contexts_rd_data          )  //o
  );
  always @(*) begin
    _zz_wr_en = 1'b0;
    if(write_valid) begin
      _zz_wr_en = 1'b1;
    end
  end

  assign write_valid = io_add_valid;
  assign write_payload_address = io_add_payload_id;
  assign write_payload_data = io_add_payload_context;
  assign io_add_ready = 1'b1;
  assign read_data = contexts_rd_data;
  assign read_address = io_query_id;
  assign io_query_context = read_data;
  assign contexts_wr_en = (_zz_wr_en && 1'b1);
  assign contexts_wr_data = write_payload_data;

endmodule

module StreamArbiter_8 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_opcode,
  input  wire [2:0]    io_inputs_0_payload_param,
  input  wire [1:0]    io_inputs_0_payload_source,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire          io_inputs_0_payload_denied,
  input  wire [63:0]   io_inputs_0_payload_data,
  input  wire          io_inputs_0_payload_corrupt,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_opcode,
  input  wire [2:0]    io_inputs_1_payload_param,
  input  wire [1:0]    io_inputs_1_payload_source,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire          io_inputs_1_payload_denied,
  input  wire [63:0]   io_inputs_1_payload_data,
  input  wire          io_inputs_1_payload_corrupt,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_opcode,
  output wire [2:0]    io_output_payload_param,
  output wire [1:0]    io_output_payload_source,
  output wire [2:0]    io_output_payload_size,
  output wire          io_output_payload_denied,
  output wire [63:0]   io_output_payload_data,
  output wire          io_output_payload_corrupt,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);
  localparam D_ACCESS_ACK = 3'd0;
  localparam D_ACCESS_ACK_DATA = 3'd1;
  localparam D_GRANT = 3'd4;
  localparam D_GRANT_DATA = 3'd5;
  localparam D_RELEASE_ACK = 3'd6;

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg        [2:0]    _zz_io_output_tracker_last;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  reg        [2:0]    io_output_tracker_beat;
  wire                io_output_tracker_last;
  wire                when_Stream_l800;
  wire       [2:0]    _zz_io_output_payload_opcode;
  wire                _zz_io_chosen;
  `ifndef SYNTHESIS
  reg [119:0] io_inputs_0_payload_opcode_string;
  reg [119:0] io_inputs_1_payload_opcode_string;
  reg [119:0] io_output_payload_opcode_string;
  reg [119:0] _zz_io_output_payload_opcode_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(io_output_payload_size)
      3'b000 : _zz_io_output_tracker_last = 3'b000;
      3'b001 : _zz_io_output_tracker_last = 3'b000;
      3'b010 : _zz_io_output_tracker_last = 3'b000;
      3'b011 : _zz_io_output_tracker_last = 3'b000;
      3'b100 : _zz_io_output_tracker_last = 3'b001;
      3'b101 : _zz_io_output_tracker_last = 3'b011;
      default : _zz_io_output_tracker_last = 3'b111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_opcode)
      D_ACCESS_ACK : io_inputs_0_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_inputs_0_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_inputs_0_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_inputs_0_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_inputs_0_payload_opcode_string = "RELEASE_ACK    ";
      default : io_inputs_0_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_opcode)
      D_ACCESS_ACK : io_inputs_1_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_inputs_1_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_inputs_1_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_inputs_1_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_inputs_1_payload_opcode_string = "RELEASE_ACK    ";
      default : io_inputs_1_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_opcode)
      D_ACCESS_ACK : io_output_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : io_output_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : io_output_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : io_output_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : io_output_payload_opcode_string = "RELEASE_ACK    ";
      default : io_output_payload_opcode_string = "???????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_opcode)
      D_ACCESS_ACK : _zz_io_output_payload_opcode_string = "ACCESS_ACK     ";
      D_ACCESS_ACK_DATA : _zz_io_output_payload_opcode_string = "ACCESS_ACK_DATA";
      D_GRANT : _zz_io_output_payload_opcode_string = "GRANT          ";
      D_GRANT_DATA : _zz_io_output_payload_opcode_string = "GRANT_DATA     ";
      D_RELEASE_ACK : _zz_io_output_payload_opcode_string = "RELEASE_ACK    ";
      default : _zz_io_output_payload_opcode_string = "???????????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_tracker_last = ((! ((1'b0 || (D_ACCESS_ACK_DATA == io_output_payload_opcode)) || (D_GRANT_DATA == io_output_payload_opcode))) || (io_output_tracker_beat == _zz_io_output_tracker_last));
  assign when_Stream_l800 = (io_output_fire && io_output_tracker_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign _zz_io_output_payload_opcode = (maskRouted_0 ? io_inputs_0_payload_opcode : io_inputs_1_payload_opcode);
  assign io_output_payload_opcode = _zz_io_output_payload_opcode;
  assign io_output_payload_param = (maskRouted_0 ? io_inputs_0_payload_param : io_inputs_1_payload_param);
  assign io_output_payload_source = (maskRouted_0 ? io_inputs_0_payload_source : io_inputs_1_payload_source);
  assign io_output_payload_size = (maskRouted_0 ? io_inputs_0_payload_size : io_inputs_1_payload_size);
  assign io_output_payload_denied = (maskRouted_0 ? io_inputs_0_payload_denied : io_inputs_1_payload_denied);
  assign io_output_payload_data = (maskRouted_0 ? io_inputs_0_payload_data : io_inputs_1_payload_data);
  assign io_output_payload_corrupt = (maskRouted_0 ? io_inputs_0_payload_corrupt : io_inputs_1_payload_corrupt);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
      io_output_tracker_beat <= 3'b000;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        io_output_tracker_beat <= (io_output_tracker_beat + 3'b001);
        if(io_output_tracker_last) begin
          io_output_tracker_beat <= 3'b000;
        end
      end
      if(when_Stream_l800) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_7 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [1:0]    io_inputs_0_payload_source,
  input  wire          io_inputs_0_payload_denied,
  input  wire          io_inputs_0_payload_last,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [1:0]    io_inputs_1_payload_source,
  input  wire          io_inputs_1_payload_denied,
  input  wire          io_inputs_1_payload_last,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [1:0]    io_output_payload_source,
  output wire          io_output_payload_denied,
  output wire          io_output_payload_last,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                when_Stream_l800;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_Stream_l800 = (io_output_fire && io_output_payload_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_source = (maskRouted_0 ? io_inputs_0_payload_source : io_inputs_1_payload_source);
  assign io_output_payload_denied = (maskRouted_0 ? io_inputs_0_payload_denied : io_inputs_1_payload_denied);
  assign io_output_payload_last = (maskRouted_0 ? io_inputs_0_payload_last : io_inputs_1_payload_last);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(when_Stream_l800) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module ContextAsyncBufferFull (
  input  wire          io_add_valid,
  output wire          io_add_ready,
  input  wire [1:0]    io_add_payload_id,
  input  wire [2:0]    io_add_payload_context,
  input  wire          io_remove_valid,
  input  wire [1:0]    io_remove_payload_id,
  input  wire [1:0]    io_query_id,
  output wire [2:0]    io_query_context,
  input  wire          litex_clk
);

  wire                contexts_wr_en;
  wire       [2:0]    contexts_wr_data;
  wire       [2:0]    contexts_rd_data;
  reg                 _zz_wr_en;
  wire                write_valid;
  wire       [1:0]    write_payload_address;
  wire       [2:0]    write_payload_data;
  wire       [1:0]    read_address;
  wire       [2:0]    read_data;

  Ram_1w_1ra #(
    .wordCount      (4         ),
    .wordWidth      (3         ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (2         ),
    .wrDataWidth    (3         ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (2         ),
    .rdDataWidth    (3         )
  ) contexts (
    .clk     (litex_clk                 ), //i
    .wr_en   (contexts_wr_en            ), //i
    .wr_mask (1'b1                      ), //i
    .wr_addr (write_payload_address[1:0]), //i
    .wr_data (contexts_wr_data[2:0]     ), //i
    .rd_addr (read_address[1:0]         ), //i
    .rd_data (contexts_rd_data[2:0]     )  //o
  );
  always @(*) begin
    _zz_wr_en = 1'b0;
    if(write_valid) begin
      _zz_wr_en = 1'b1;
    end
  end

  assign write_valid = io_add_valid;
  assign write_payload_address = io_add_payload_id;
  assign write_payload_data = io_add_payload_context;
  assign io_add_ready = 1'b1;
  assign read_data = contexts_rd_data;
  assign read_address = io_query_id;
  assign io_query_context = read_data;
  assign contexts_wr_en = (_zz_wr_en && 1'b1);
  assign contexts_wr_data = write_payload_data;

endmodule

module StreamArbiter_6 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_opcode,
  input  wire [2:0]    io_inputs_0_payload_param,
  input  wire [2:0]    io_inputs_0_payload_source,
  input  wire [31:0]   io_inputs_0_payload_address,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire [3:0]    io_inputs_0_payload_mask,
  input  wire [31:0]   io_inputs_0_payload_data,
  input  wire          io_inputs_0_payload_corrupt,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_opcode,
  input  wire [2:0]    io_inputs_1_payload_param,
  input  wire [2:0]    io_inputs_1_payload_source,
  input  wire [31:0]   io_inputs_1_payload_address,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire [3:0]    io_inputs_1_payload_mask,
  input  wire [31:0]   io_inputs_1_payload_data,
  input  wire          io_inputs_1_payload_corrupt,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_opcode,
  output wire [2:0]    io_output_payload_param,
  output wire [2:0]    io_output_payload_source,
  output wire [31:0]   io_output_payload_address,
  output wire [2:0]    io_output_payload_size,
  output wire [3:0]    io_output_payload_mask,
  output wire [31:0]   io_output_payload_data,
  output wire          io_output_payload_corrupt,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          litex_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg        [3:0]    _zz_io_output_tracker_last;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  reg        [3:0]    io_output_tracker_beat;
  wire                io_output_tracker_last;
  wire                when_Stream_l800;
  wire       [2:0]    _zz_io_output_payload_opcode;
  wire                _zz_io_chosen;
  `ifndef SYNTHESIS
  reg [127:0] io_inputs_0_payload_opcode_string;
  reg [127:0] io_inputs_1_payload_opcode_string;
  reg [127:0] io_output_payload_opcode_string;
  reg [127:0] _zz_io_output_payload_opcode_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(io_output_payload_size)
      3'b000 : _zz_io_output_tracker_last = 4'b0000;
      3'b001 : _zz_io_output_tracker_last = 4'b0000;
      3'b010 : _zz_io_output_tracker_last = 4'b0000;
      3'b011 : _zz_io_output_tracker_last = 4'b0001;
      3'b100 : _zz_io_output_tracker_last = 4'b0011;
      3'b101 : _zz_io_output_tracker_last = 4'b0111;
      default : _zz_io_output_tracker_last = 4'b1111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_opcode)
      A_PUT_FULL_DATA : io_inputs_0_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_inputs_0_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_inputs_0_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_inputs_0_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_inputs_0_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_inputs_0_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_opcode)
      A_PUT_FULL_DATA : io_inputs_1_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_inputs_1_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_inputs_1_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_inputs_1_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_inputs_1_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_inputs_1_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_opcode)
      A_PUT_FULL_DATA : io_output_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_output_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_output_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_output_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_output_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_output_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_opcode)
      A_PUT_FULL_DATA : _zz_io_output_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_output_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_output_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_output_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_output_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_io_output_payload_opcode_string = "????????????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == io_output_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_output_payload_opcode))) || (io_output_tracker_beat == _zz_io_output_tracker_last));
  assign when_Stream_l800 = (io_output_fire && io_output_tracker_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign _zz_io_output_payload_opcode = (maskRouted_0 ? io_inputs_0_payload_opcode : io_inputs_1_payload_opcode);
  assign io_output_payload_opcode = _zz_io_output_payload_opcode;
  assign io_output_payload_param = (maskRouted_0 ? io_inputs_0_payload_param : io_inputs_1_payload_param);
  assign io_output_payload_source = (maskRouted_0 ? io_inputs_0_payload_source : io_inputs_1_payload_source);
  assign io_output_payload_address = (maskRouted_0 ? io_inputs_0_payload_address : io_inputs_1_payload_address);
  assign io_output_payload_size = (maskRouted_0 ? io_inputs_0_payload_size : io_inputs_1_payload_size);
  assign io_output_payload_mask = (maskRouted_0 ? io_inputs_0_payload_mask : io_inputs_1_payload_mask);
  assign io_output_payload_data = (maskRouted_0 ? io_inputs_0_payload_data : io_inputs_1_payload_data);
  assign io_output_payload_corrupt = (maskRouted_0 ? io_inputs_0_payload_corrupt : io_inputs_1_payload_corrupt);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge litex_clk or posedge litex_reset) begin
    if(litex_reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
      io_output_tracker_beat <= 4'b0000;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        io_output_tracker_beat <= (io_output_tracker_beat + 4'b0001);
        if(io_output_tracker_last) begin
          io_output_tracker_beat <= 4'b0000;
        end
      end
      if(when_Stream_l800) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_5 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_opcode,
  input  wire [2:0]    io_inputs_0_payload_param,
  input  wire [1:0]    io_inputs_0_payload_source,
  input  wire [31:0]   io_inputs_0_payload_address,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire [7:0]    io_inputs_0_payload_mask,
  input  wire [63:0]   io_inputs_0_payload_data,
  input  wire          io_inputs_0_payload_corrupt,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_opcode,
  input  wire [2:0]    io_inputs_1_payload_param,
  input  wire [1:0]    io_inputs_1_payload_source,
  input  wire [31:0]   io_inputs_1_payload_address,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire [7:0]    io_inputs_1_payload_mask,
  input  wire [63:0]   io_inputs_1_payload_data,
  input  wire          io_inputs_1_payload_corrupt,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_opcode,
  output wire [2:0]    io_output_payload_param,
  output wire [1:0]    io_output_payload_source,
  output wire [31:0]   io_output_payload_address,
  output wire [2:0]    io_output_payload_size,
  output wire [7:0]    io_output_payload_mask,
  output wire [63:0]   io_output_payload_data,
  output wire          io_output_payload_corrupt,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);
  localparam A_PUT_FULL_DATA = 3'd0;
  localparam A_PUT_PARTIAL_DATA = 3'd1;
  localparam A_GET = 3'd4;
  localparam A_ACQUIRE_BLOCK = 3'd6;
  localparam A_ACQUIRE_PERM = 3'd7;

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg        [2:0]    _zz_io_output_tracker_last;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  reg        [2:0]    io_output_tracker_beat;
  wire                io_output_tracker_last;
  wire                when_Stream_l800;
  wire       [2:0]    _zz_io_output_payload_opcode;
  wire                _zz_io_chosen;
  `ifndef SYNTHESIS
  reg [127:0] io_inputs_0_payload_opcode_string;
  reg [127:0] io_inputs_1_payload_opcode_string;
  reg [127:0] io_output_payload_opcode_string;
  reg [127:0] _zz_io_output_payload_opcode_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(io_output_payload_size)
      3'b000 : _zz_io_output_tracker_last = 3'b000;
      3'b001 : _zz_io_output_tracker_last = 3'b000;
      3'b010 : _zz_io_output_tracker_last = 3'b000;
      3'b011 : _zz_io_output_tracker_last = 3'b000;
      3'b100 : _zz_io_output_tracker_last = 3'b001;
      3'b101 : _zz_io_output_tracker_last = 3'b011;
      default : _zz_io_output_tracker_last = 3'b111;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_opcode)
      A_PUT_FULL_DATA : io_inputs_0_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_inputs_0_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_inputs_0_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_inputs_0_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_inputs_0_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_inputs_0_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_opcode)
      A_PUT_FULL_DATA : io_inputs_1_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_inputs_1_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_inputs_1_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_inputs_1_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_inputs_1_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_inputs_1_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_opcode)
      A_PUT_FULL_DATA : io_output_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : io_output_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : io_output_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : io_output_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : io_output_payload_opcode_string = "ACQUIRE_PERM    ";
      default : io_output_payload_opcode_string = "????????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_opcode)
      A_PUT_FULL_DATA : _zz_io_output_payload_opcode_string = "PUT_FULL_DATA   ";
      A_PUT_PARTIAL_DATA : _zz_io_output_payload_opcode_string = "PUT_PARTIAL_DATA";
      A_GET : _zz_io_output_payload_opcode_string = "GET             ";
      A_ACQUIRE_BLOCK : _zz_io_output_payload_opcode_string = "ACQUIRE_BLOCK   ";
      A_ACQUIRE_PERM : _zz_io_output_payload_opcode_string = "ACQUIRE_PERM    ";
      default : _zz_io_output_payload_opcode_string = "????????????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_tracker_last = ((! ((1'b0 || (A_PUT_FULL_DATA == io_output_payload_opcode)) || (A_PUT_PARTIAL_DATA == io_output_payload_opcode))) || (io_output_tracker_beat == _zz_io_output_tracker_last));
  assign when_Stream_l800 = (io_output_fire && io_output_tracker_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign _zz_io_output_payload_opcode = (maskRouted_0 ? io_inputs_0_payload_opcode : io_inputs_1_payload_opcode);
  assign io_output_payload_opcode = _zz_io_output_payload_opcode;
  assign io_output_payload_param = (maskRouted_0 ? io_inputs_0_payload_param : io_inputs_1_payload_param);
  assign io_output_payload_source = (maskRouted_0 ? io_inputs_0_payload_source : io_inputs_1_payload_source);
  assign io_output_payload_address = (maskRouted_0 ? io_inputs_0_payload_address : io_inputs_1_payload_address);
  assign io_output_payload_size = (maskRouted_0 ? io_inputs_0_payload_size : io_inputs_1_payload_size);
  assign io_output_payload_mask = (maskRouted_0 ? io_inputs_0_payload_mask : io_inputs_1_payload_mask);
  assign io_output_payload_data = (maskRouted_0 ? io_inputs_0_payload_data : io_inputs_1_payload_data);
  assign io_output_payload_corrupt = (maskRouted_0 ? io_inputs_0_payload_corrupt : io_inputs_1_payload_corrupt);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
      io_output_tracker_beat <= 3'b000;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        io_output_tracker_beat <= (io_output_tracker_beat + 3'b001);
        if(io_output_tracker_last) begin
          io_output_tracker_beat <= 3'b000;
        end
      end
      if(when_Stream_l800) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module RegFileMem (
  input  wire          io_writes_0_valid,
  input  wire [4:0]    io_writes_0_address,
  input  wire [31:0]   io_writes_0_data,
  input  wire [15:0]   io_writes_0_uopId,
  input  wire          io_reads_0_valid,
  input  wire [4:0]    io_reads_0_address,
  output wire [31:0]   io_reads_0_data,
  input  wire          io_reads_1_valid,
  input  wire [4:0]    io_reads_1_address,
  output wire [31:0]   io_reads_1_data,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);

  reg        [31:0]   asMem_ram_spinal_port1;
  reg        [31:0]   asMem_ram_spinal_port2;
  reg                 _zz_1;
  wire                conv_writes_0_valid;
  wire       [4:0]    conv_writes_0_payload_address;
  wire       [31:0]   conv_writes_0_payload_data;
  wire                conv_read_0_cmd_valid;
  wire       [4:0]    conv_read_0_cmd_payload;
  wire       [31:0]   conv_read_0_rsp;
  wire                conv_read_1_cmd_valid;
  wire       [4:0]    conv_read_1_cmd_payload;
  wire       [31:0]   conv_read_1_rsp;
  wire                asMem_writes_0_port_valid;
  wire       [4:0]    asMem_writes_0_port_payload_address;
  wire       [31:0]   asMem_writes_0_port_payload_data;
  wire                asMem_reads_0_sync_port_cmd_valid;
  wire       [4:0]    asMem_reads_0_sync_port_cmd_payload;
  wire       [31:0]   asMem_reads_0_sync_port_rsp;
  wire                asMem_reads_1_sync_port_cmd_valid;
  wire       [4:0]    asMem_reads_1_sync_port_cmd_payload;
  wire       [31:0]   asMem_reads_1_sync_port_rsp;
  reg [31:0] asMem_ram [0:31] /* verilator public */ ;

  always @(posedge litex_clk) begin
    if(_zz_1) begin
      asMem_ram[asMem_writes_0_port_payload_address] <= asMem_writes_0_port_payload_data;
    end
  end

  always @(posedge litex_clk) begin
    if(asMem_reads_0_sync_port_cmd_valid) begin
      asMem_ram_spinal_port1 <= asMem_ram[asMem_reads_0_sync_port_cmd_payload];
    end
  end

  always @(posedge litex_clk) begin
    if(asMem_reads_1_sync_port_cmd_valid) begin
      asMem_ram_spinal_port2 <= asMem_ram[asMem_reads_1_sync_port_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(asMem_writes_0_port_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign conv_writes_0_valid = io_writes_0_valid;
  assign conv_writes_0_payload_address = io_writes_0_address;
  assign conv_writes_0_payload_data = io_writes_0_data;
  assign conv_read_0_cmd_valid = io_reads_0_valid;
  assign conv_read_0_cmd_payload = io_reads_0_address;
  assign io_reads_0_data = conv_read_0_rsp;
  assign conv_read_1_cmd_valid = io_reads_1_valid;
  assign conv_read_1_cmd_payload = io_reads_1_address;
  assign io_reads_1_data = conv_read_1_rsp;
  assign asMem_writes_0_port_valid = conv_writes_0_valid;
  assign asMem_writes_0_port_payload_address = conv_writes_0_payload_address;
  assign asMem_writes_0_port_payload_data = conv_writes_0_payload_data;
  assign asMem_reads_0_sync_port_rsp = asMem_ram_spinal_port1;
  assign asMem_reads_0_sync_port_cmd_valid = conv_read_0_cmd_valid;
  assign asMem_reads_0_sync_port_cmd_payload = conv_read_0_cmd_payload;
  assign conv_read_0_rsp = asMem_reads_0_sync_port_rsp;
  assign asMem_reads_1_sync_port_rsp = asMem_ram_spinal_port2;
  assign asMem_reads_1_sync_port_cmd_valid = conv_read_1_cmd_valid;
  assign asMem_reads_1_sync_port_cmd_payload = conv_read_1_cmd_payload;
  assign conv_read_1_rsp = asMem_reads_1_sync_port_rsp;

endmodule

module StreamArbiter_4 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [0:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;
  wire                io_output_fire;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_3 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [31:0]   io_inputs_0_payload_address,
  input  wire [0:0]    io_inputs_0_payload_storageId,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [31:0]   io_output_payload_address,
  output wire [0:0]    io_output_payload_storageId,
  output wire [0:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;
  wire                io_output_fire;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_output_payload_address = io_inputs_0_payload_address;
  assign io_output_payload_storageId = io_inputs_0_payload_storageId;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_2 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [2:0]    io_inputs_0_payload_op,
  input  wire [31:0]   io_inputs_0_payload_address,
  input  wire [1:0]    io_inputs_0_payload_size,
  input  wire          io_inputs_0_payload_load,
  input  wire          io_inputs_0_payload_store,
  input  wire          io_inputs_0_payload_atomic,
  input  wire          io_inputs_0_payload_clean,
  input  wire          io_inputs_0_payload_invalidate,
  input  wire [11:0]   io_inputs_0_payload_storeId,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [2:0]    io_inputs_1_payload_op,
  input  wire [31:0]   io_inputs_1_payload_address,
  input  wire [1:0]    io_inputs_1_payload_size,
  input  wire          io_inputs_1_payload_load,
  input  wire          io_inputs_1_payload_store,
  input  wire          io_inputs_1_payload_atomic,
  input  wire          io_inputs_1_payload_clean,
  input  wire          io_inputs_1_payload_invalidate,
  input  wire [11:0]   io_inputs_1_payload_storeId,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [2:0]    io_inputs_2_payload_op,
  input  wire [31:0]   io_inputs_2_payload_address,
  input  wire [1:0]    io_inputs_2_payload_size,
  input  wire          io_inputs_2_payload_load,
  input  wire          io_inputs_2_payload_store,
  input  wire          io_inputs_2_payload_atomic,
  input  wire          io_inputs_2_payload_clean,
  input  wire          io_inputs_2_payload_invalidate,
  input  wire [11:0]   io_inputs_2_payload_storeId,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [2:0]    io_output_payload_op,
  output wire [31:0]   io_output_payload_address,
  output wire [1:0]    io_output_payload_size,
  output wire          io_output_payload_load,
  output wire          io_output_payload_store,
  output wire          io_output_payload_atomic,
  output wire          io_output_payload_clean,
  output wire          io_output_payload_invalidate,
  output wire [11:0]   io_output_payload_storeId,
  output wire [1:0]    io_chosen,
  output wire [2:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);
  localparam LsuL1CmdOpcode_LSU = 3'd0;
  localparam LsuL1CmdOpcode_ACCESS_1 = 3'd1;
  localparam LsuL1CmdOpcode_STORE_BUFFER = 3'd2;
  localparam LsuL1CmdOpcode_FLUSH = 3'd3;
  localparam LsuL1CmdOpcode_PREFETCH = 3'd4;

  wire       [2:0]    _zz__zz_maskProposal_1_1;
  reg        [2:0]    _zz__zz_io_output_payload_op;
  reg        [31:0]   _zz_io_output_payload_address_1;
  reg        [1:0]    _zz_io_output_payload_size;
  reg                 _zz_io_output_payload_load;
  reg                 _zz_io_output_payload_store;
  reg                 _zz_io_output_payload_atomic;
  reg                 _zz_io_output_payload_clean;
  reg                 _zz_io_output_payload_invalidate;
  reg        [11:0]   _zz_io_output_payload_storeId;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire       [2:0]    _zz_maskProposal_1;
  wire       [2:0]    _zz_maskProposal_1_1;
  wire       [1:0]    _zz_io_output_payload_address;
  wire       [2:0]    _zz_io_output_payload_op;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  `ifndef SYNTHESIS
  reg [95:0] io_inputs_0_payload_op_string;
  reg [95:0] io_inputs_1_payload_op_string;
  reg [95:0] io_inputs_2_payload_op_string;
  reg [95:0] io_output_payload_op_string;
  reg [95:0] _zz_io_output_payload_op_string;
  `endif


  assign _zz__zz_maskProposal_1_1 = (_zz_maskProposal_1 - 3'b001);
  always @(*) begin
    case(_zz_io_output_payload_address)
      2'b00 : begin
        _zz__zz_io_output_payload_op = io_inputs_0_payload_op;
        _zz_io_output_payload_address_1 = io_inputs_0_payload_address;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_load = io_inputs_0_payload_load;
        _zz_io_output_payload_store = io_inputs_0_payload_store;
        _zz_io_output_payload_atomic = io_inputs_0_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_0_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_0_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_0_payload_storeId;
      end
      2'b01 : begin
        _zz__zz_io_output_payload_op = io_inputs_1_payload_op;
        _zz_io_output_payload_address_1 = io_inputs_1_payload_address;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_load = io_inputs_1_payload_load;
        _zz_io_output_payload_store = io_inputs_1_payload_store;
        _zz_io_output_payload_atomic = io_inputs_1_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_1_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_1_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_1_payload_storeId;
      end
      default : begin
        _zz__zz_io_output_payload_op = io_inputs_2_payload_op;
        _zz_io_output_payload_address_1 = io_inputs_2_payload_address;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_load = io_inputs_2_payload_load;
        _zz_io_output_payload_store = io_inputs_2_payload_store;
        _zz_io_output_payload_atomic = io_inputs_2_payload_atomic;
        _zz_io_output_payload_clean = io_inputs_2_payload_clean;
        _zz_io_output_payload_invalidate = io_inputs_2_payload_invalidate;
        _zz_io_output_payload_storeId = io_inputs_2_payload_storeId;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_0_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_0_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_0_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_0_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_0_payload_op_string = "PREFETCH    ";
      default : io_inputs_0_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_1_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_1_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_1_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_1_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_1_payload_op_string = "PREFETCH    ";
      default : io_inputs_1_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_op)
      LsuL1CmdOpcode_LSU : io_inputs_2_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_inputs_2_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_inputs_2_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_inputs_2_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_inputs_2_payload_op_string = "PREFETCH    ";
      default : io_inputs_2_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_op)
      LsuL1CmdOpcode_LSU : io_output_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : io_output_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : io_output_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : io_output_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : io_output_payload_op_string = "PREFETCH    ";
      default : io_output_payload_op_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_op)
      LsuL1CmdOpcode_LSU : _zz_io_output_payload_op_string = "LSU         ";
      LsuL1CmdOpcode_ACCESS_1 : _zz_io_output_payload_op_string = "ACCESS_1    ";
      LsuL1CmdOpcode_STORE_BUFFER : _zz_io_output_payload_op_string = "STORE_BUFFER";
      LsuL1CmdOpcode_FLUSH : _zz_io_output_payload_op_string = "FLUSH       ";
      LsuL1CmdOpcode_PREFETCH : _zz_io_output_payload_op_string = "PREFETCH    ";
      default : _zz_io_output_payload_op_string = "????????????";
    endcase
  end
  `endif

  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign _zz_maskProposal_1 = {io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}};
  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz__zz_maskProposal_1_1));
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign maskProposal_2 = _zz_maskProposal_1_1[2];
  assign io_output_valid = (((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2));
  assign _zz_io_output_payload_address = {maskRouted_2,maskRouted_1};
  assign _zz_io_output_payload_op = _zz__zz_io_output_payload_op;
  assign io_output_payload_op = _zz_io_output_payload_op;
  assign io_output_payload_address = _zz_io_output_payload_address_1;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_load = _zz_io_output_payload_load;
  assign io_output_payload_store = _zz_io_output_payload_store;
  assign io_output_payload_atomic = _zz_io_output_payload_atomic;
  assign io_output_payload_clean = _zz_io_output_payload_clean;
  assign io_output_payload_invalidate = _zz_io_output_payload_invalidate;
  assign io_output_payload_storeId = _zz_io_output_payload_storeId;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_chosenOH = {maskRouted_2,{maskRouted_1,maskRouted_0}};
  assign _zz_io_chosen = io_chosenOH[1];
  assign _zz_io_chosen_1 = io_chosenOH[2];
  assign io_chosen = {_zz_io_chosen_1,_zz_io_chosen};
  always @(posedge litex_clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
      maskLocked_2 <= maskRouted_2;
    end
  end


endmodule

module StreamArbiter_1 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [31:0]   io_inputs_0_payload_pcOnLastSlice,
  input  wire [31:0]   io_inputs_0_payload_pcTarget,
  input  wire          io_inputs_0_payload_taken,
  input  wire          io_inputs_0_payload_isBranch,
  input  wire          io_inputs_0_payload_isPush,
  input  wire          io_inputs_0_payload_isPop,
  input  wire          io_inputs_0_payload_wasWrong,
  input  wire          io_inputs_0_payload_badPredictedTarget,
  input  wire [11:0]   io_inputs_0_payload_history,
  input  wire [15:0]   io_inputs_0_payload_uopId,
  input  wire [1:0]    io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [31:0]   io_output_payload_pcOnLastSlice,
  output wire [31:0]   io_output_payload_pcTarget,
  output wire          io_output_payload_taken,
  output wire          io_output_payload_isBranch,
  output wire          io_output_payload_isPush,
  output wire          io_output_payload_isPop,
  output wire          io_output_payload_wasWrong,
  output wire          io_output_payload_badPredictedTarget,
  output wire [11:0]   io_output_payload_history,
  output wire [15:0]   io_output_payload_uopId,
  output wire [1:0]    io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0,
  output wire [0:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  wire                locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_output_payload_pcOnLastSlice = io_inputs_0_payload_pcOnLastSlice;
  assign io_output_payload_pcTarget = io_inputs_0_payload_pcTarget;
  assign io_output_payload_taken = io_inputs_0_payload_taken;
  assign io_output_payload_isBranch = io_inputs_0_payload_isBranch;
  assign io_output_payload_isPush = io_inputs_0_payload_isPush;
  assign io_output_payload_isPop = io_inputs_0_payload_isPop;
  assign io_output_payload_wasWrong = io_inputs_0_payload_wasWrong;
  assign io_output_payload_badPredictedTarget = io_inputs_0_payload_badPredictedTarget;
  assign io_output_payload_history = io_inputs_0_payload_history;
  assign io_output_payload_uopId = io_inputs_0_payload_uopId;
  assign io_output_payload_ctx_GSharePlugin_GSHARE_COUNTER_0 = io_inputs_0_payload_ctx_GSharePlugin_GSHARE_COUNTER_0;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
    end
  end


endmodule

module StreamArbiter (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [0:0]    io_chosenOH,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);

  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire                io_output_fire;

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskProposal_0 = io_inputs_0_valid;
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      locked <= 1'b0;
    end else begin
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end

  always @(posedge litex_clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
    end
  end


endmodule

module StreamFifoLowLatency (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_outputs_0,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_outputs_0,
  input  wire          io_flush,
  output wire [1:0]    io_occupancy,
  output wire [1:0]    io_availability,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);

  wire                fifo_io_push_ready;
  wire                fifo_io_pop_valid;
  wire       [31:0]   fifo_io_pop_payload_outputs_0;
  wire       [1:0]    fifo_io_occupancy;
  wire       [1:0]    fifo_io_availability;

  StreamFifo fifo (
    .io_push_valid             (io_push_valid                      ), //i
    .io_push_ready             (fifo_io_push_ready                 ), //o
    .io_push_payload_outputs_0 (io_push_payload_outputs_0[31:0]    ), //i
    .io_pop_valid              (fifo_io_pop_valid                  ), //o
    .io_pop_ready              (io_pop_ready                       ), //i
    .io_pop_payload_outputs_0  (fifo_io_pop_payload_outputs_0[31:0]), //o
    .io_flush                  (io_flush                           ), //i
    .io_occupancy              (fifo_io_occupancy[1:0]             ), //o
    .io_availability           (fifo_io_availability[1:0]          ), //o
    .litex_clk                 (litex_clk                          ), //i
    .cpuResetCtrl_reset        (cpuResetCtrl_reset                 )  //i
  );
  assign io_push_ready = fifo_io_push_ready;
  assign io_pop_valid = fifo_io_pop_valid;
  assign io_pop_payload_outputs_0 = fifo_io_pop_payload_outputs_0;
  assign io_occupancy = fifo_io_occupancy;
  assign io_availability = fifo_io_availability;

endmodule

module DivRadix (
  input  wire          io_flush,
  input  wire          io_cmd_valid,
  output wire          io_cmd_ready,
  input  wire [31:0]   io_cmd_payload_a,
  input  wire [31:0]   io_cmd_payload_b,
  input  wire          io_cmd_payload_normalized,
  input  wire [4:0]    io_cmd_payload_iterations,
  output wire          io_rsp_valid,
  input  wire          io_rsp_ready,
  output wire [31:0]   io_rsp_payload_result,
  output wire [31:0]   io_rsp_payload_remain,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);

  wire       [7:0]    _zz_shifter_1;
  wire       [15:0]   _zz_shifter_2;
  wire       [23:0]   _zz_shifter_3;
  wire       [30:0]   _zz_shifter_4;
  reg        [4:0]    counter;
  reg                 busy;
  wire                io_rsp_fire;
  reg                 done;
  wire                when_DivRadix_l45;
  reg        [31:0]   shifter;
  reg        [31:0]   numerator;
  reg        [31:0]   result;
  reg        [32:0]   div1;
  reg        [32:0]   div3;
  wire       [32:0]   div2;
  wire       [32:0]   shifted;
  wire       [33:0]   sub1;
  wire                when_DivRadix_l64;
  reg        [32:0]   _zz_shifter;
  wire                when_DivRadix_l68;
  wire                slicesZero_0;
  wire                slicesZero_1;
  wire                slicesZero_2;
  wire       [2:0]    shiftSel;
  wire       [3:0]    _zz_sel;
  wire                _zz_sel_1;
  wire                _zz_sel_2;
  wire                _zz_sel_3;
  reg        [3:0]    _zz_sel_4;
  wire       [3:0]    _zz_sel_5;
  wire                _zz_sel_6;
  wire                _zz_sel_7;
  wire                _zz_sel_8;
  wire       [1:0]    sel;
  reg                 wasBusy;
  wire                when_DivRadix_l93;

  assign _zz_shifter_1 = io_cmd_payload_a[31 : 24];
  assign _zz_shifter_2 = io_cmd_payload_a[31 : 16];
  assign _zz_shifter_3 = io_cmd_payload_a[31 : 8];
  assign _zz_shifter_4 = io_cmd_payload_a[31 : 1];
  assign io_rsp_fire = (io_rsp_valid && io_rsp_ready);
  assign when_DivRadix_l45 = (busy && (counter == 5'h1f));
  assign div2 = (div1 <<< 1);
  assign shifted = {shifter,numerator[31 : 31]};
  assign sub1 = ({1'b0,shifted} - {1'b0,div1});
  assign io_rsp_valid = done;
  assign io_rsp_payload_result = result;
  assign io_rsp_payload_remain = shifter;
  assign io_cmd_ready = (! busy);
  assign when_DivRadix_l64 = (! done);
  always @(*) begin
    _zz_shifter = shifted;
    if(when_DivRadix_l68) begin
      _zz_shifter = sub1[32:0];
    end
  end

  assign when_DivRadix_l68 = (! sub1[33]);
  assign slicesZero_0 = (io_cmd_payload_a[15 : 8] == 8'h0);
  assign slicesZero_1 = (io_cmd_payload_a[23 : 16] == 8'h0);
  assign slicesZero_2 = (io_cmd_payload_a[31 : 24] == 8'h0);
  assign shiftSel = {(&slicesZero_2),{(&{slicesZero_2,slicesZero_1}),(&{slicesZero_2,{slicesZero_1,slicesZero_0}})}};
  assign _zz_sel = {1'b1,shiftSel};
  assign _zz_sel_1 = _zz_sel[0];
  assign _zz_sel_2 = _zz_sel[1];
  assign _zz_sel_3 = _zz_sel[2];
  always @(*) begin
    _zz_sel_4[0] = (_zz_sel_1 && (! 1'b0));
    _zz_sel_4[1] = (_zz_sel_2 && (! _zz_sel_1));
    _zz_sel_4[2] = (_zz_sel_3 && (! (|{_zz_sel_2,_zz_sel_1})));
    _zz_sel_4[3] = (_zz_sel[3] && (! (|{_zz_sel_3,{_zz_sel_2,_zz_sel_1}})));
  end

  assign _zz_sel_5 = _zz_sel_4;
  assign _zz_sel_6 = _zz_sel_5[3];
  assign _zz_sel_7 = (_zz_sel_5[1] || _zz_sel_6);
  assign _zz_sel_8 = (_zz_sel_5[2] || _zz_sel_6);
  assign sel = {_zz_sel_8,_zz_sel_7};
  assign when_DivRadix_l93 = (! busy);
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      busy <= 1'b0;
      done <= 1'b0;
      wasBusy <= 1'b0;
    end else begin
      if(io_rsp_fire) begin
        busy <= 1'b0;
      end
      if(when_DivRadix_l45) begin
        done <= 1'b1;
      end
      if(io_rsp_fire) begin
        done <= 1'b0;
      end
      wasBusy <= busy;
      if(when_DivRadix_l93) begin
        busy <= io_cmd_valid;
      end
      if(io_flush) begin
        done <= 1'b0;
        busy <= 1'b0;
      end
    end
  end

  always @(posedge litex_clk) begin
    if(when_DivRadix_l64) begin
      counter <= (counter + 5'h01);
      result <= (result <<< 1);
      if(when_DivRadix_l68) begin
        result[0 : 0] <= 1'b1;
      end
      shifter <= _zz_shifter[31:0];
      numerator <= (numerator <<< 1);
    end
    if(when_DivRadix_l93) begin
      div1 <= {1'd0, io_cmd_payload_b};
      result <= ((io_cmd_payload_b == 32'h0) ? 32'hffffffff : 32'h0);
      case(sel)
        2'b11 : begin
          counter <= 5'h0;
          shifter <= 32'h0;
          numerator <= (io_cmd_payload_a <<< 0);
        end
        2'b10 : begin
          counter <= 5'h08;
          shifter <= {24'd0, _zz_shifter_1};
          numerator <= (io_cmd_payload_a <<< 8);
        end
        2'b01 : begin
          counter <= 5'h10;
          shifter <= {16'd0, _zz_shifter_2};
          numerator <= (io_cmd_payload_a <<< 16);
        end
        default : begin
          counter <= 5'h18;
          shifter <= {8'd0, _zz_shifter_3};
          numerator <= (io_cmd_payload_a <<< 24);
        end
      endcase
      if(io_cmd_payload_normalized) begin
        counter <= (5'h1f - io_cmd_payload_iterations);
        shifter <= {1'd0, _zz_shifter_4};
        numerator <= (io_cmd_payload_a <<< 31);
      end
    end
  end


endmodule

module StreamFifo (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_outputs_0,
  output reg           io_pop_valid,
  input  wire          io_pop_ready,
  output reg  [31:0]   io_pop_payload_outputs_0,
  input  wire          io_flush,
  output wire [1:0]    io_occupancy,
  output wire [1:0]    io_availability,
  input  wire          litex_clk,
  input  wire          cpuResetCtrl_reset
);

  wire                logic_ram_wr_en;
  wire       [31:0]   logic_ram_rd_data;
  wire       [1:0]    _zz_logic_ptr_notPow2_counter;
  wire       [1:0]    _zz_logic_ptr_notPow2_counter_1;
  wire       [0:0]    _zz_logic_ptr_notPow2_counter_2;
  wire       [1:0]    _zz_logic_ptr_notPow2_counter_3;
  wire       [0:0]    _zz_logic_ptr_notPow2_counter_4;
  wire       [31:0]   _zz_logic_pop_async_readed_outputs_0;
  reg                 _zz_wr_en;
  reg                 logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [1:0]    logic_ptr_push;
  reg        [1:0]    logic_ptr_pop;
  wire       [1:0]    logic_ptr_occupancy;
  wire       [1:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1279;
  reg                 logic_ptr_wentUp;
  wire                when_Stream_l1314;
  wire                when_Stream_l1318;
  reg        [1:0]    logic_ptr_notPow2_counter;
  wire                io_push_fire;
  wire                io_pop_fire;
  wire                logic_push_onRam_write_valid;
  wire       [1:0]    logic_push_onRam_write_payload_address;
  wire       [31:0]   logic_push_onRam_write_payload_data_outputs_0;
  wire                logic_pop_addressGen_valid;
  wire                logic_pop_addressGen_ready;
  wire       [1:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire       [31:0]   logic_pop_async_readed_outputs_0;
  wire                logic_pop_addressGen_translated_valid;
  wire                logic_pop_addressGen_translated_ready;
  wire       [31:0]   logic_pop_addressGen_translated_payload_outputs_0;

  assign _zz_logic_ptr_notPow2_counter = (logic_ptr_notPow2_counter + _zz_logic_ptr_notPow2_counter_1);
  assign _zz_logic_ptr_notPow2_counter_2 = io_push_fire;
  assign _zz_logic_ptr_notPow2_counter_1 = {1'd0, _zz_logic_ptr_notPow2_counter_2};
  assign _zz_logic_ptr_notPow2_counter_4 = io_pop_fire;
  assign _zz_logic_ptr_notPow2_counter_3 = {1'd0, _zz_logic_ptr_notPow2_counter_4};
  assign _zz_logic_pop_async_readed_outputs_0 = logic_ram_rd_data[31 : 0];
  Ram_1w_1ra #(
    .wordCount      (3         ),
    .wordWidth      (32        ),
    .technology     ("auto"    ),
    .readUnderWrite ("dontCare"),
    .wrAddressWidth (2         ),
    .wrDataWidth    (32        ),
    .wrMaskWidth    (1         ),
    .wrMaskEnable   (1'b0      ),
    .rdAddressWidth (2         ),
    .rdDataWidth    (32        )
  ) logic_ram (
    .clk     (litex_clk                                          ), //i
    .wr_en   (logic_ram_wr_en                                    ), //i
    .wr_mask (1'b1                                               ), //i
    .wr_addr (logic_push_onRam_write_payload_address[1:0]        ), //i
    .wr_data (logic_push_onRam_write_payload_data_outputs_0[31:0]), //i
    .rd_addr (logic_pop_addressGen_payload[1:0]                  ), //i
    .rd_data (logic_ram_rd_data[31:0]                            )  //o
  );
  always @(*) begin
    _zz_wr_en = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_wr_en = 1'b1;
    end
  end

  assign when_Stream_l1279 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = ((logic_ptr_push == logic_ptr_popOnIo) && logic_ptr_wentUp);
  assign logic_ptr_empty = ((logic_ptr_push == logic_ptr_pop) && (! logic_ptr_wentUp));
  assign when_Stream_l1314 = (logic_ptr_push == 2'b10);
  assign when_Stream_l1318 = (logic_ptr_pop == 2'b10);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign io_pop_fire = (io_pop_valid && io_pop_ready);
  assign logic_ptr_occupancy = logic_ptr_notPow2_counter;
  assign io_push_ready = (! logic_ptr_full);
  always @(*) begin
    logic_ptr_doPush = io_push_fire;
    if(logic_ptr_empty) begin
      if(io_pop_ready) begin
        logic_ptr_doPush = 1'b0;
      end
    end
  end

  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push;
  assign logic_push_onRam_write_payload_data_outputs_0 = io_push_payload_outputs_0;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop;
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  assign logic_pop_async_readed_outputs_0 = _zz_logic_pop_async_readed_outputs_0[31 : 0];
  assign logic_pop_addressGen_translated_valid = logic_pop_addressGen_valid;
  assign logic_pop_addressGen_ready = logic_pop_addressGen_translated_ready;
  assign logic_pop_addressGen_translated_payload_outputs_0 = logic_pop_async_readed_outputs_0;
  always @(*) begin
    io_pop_valid = logic_pop_addressGen_translated_valid;
    if(logic_ptr_empty) begin
      io_pop_valid = io_push_valid;
    end
  end

  assign logic_pop_addressGen_translated_ready = io_pop_ready;
  always @(*) begin
    io_pop_payload_outputs_0 = logic_pop_addressGen_translated_payload_outputs_0;
    if(logic_ptr_empty) begin
      io_pop_payload_outputs_0 = io_push_payload_outputs_0;
    end
  end

  assign logic_ptr_popOnIo = logic_ptr_pop;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (2'b11 - logic_ptr_occupancy);
  assign logic_ram_wr_en = (_zz_wr_en && 1'b1);
  always @(posedge litex_clk or posedge cpuResetCtrl_reset) begin
    if(cpuResetCtrl_reset) begin
      logic_ptr_push <= 2'b00;
      logic_ptr_pop <= 2'b00;
      logic_ptr_wentUp <= 1'b0;
      logic_ptr_notPow2_counter <= 2'b00;
    end else begin
      if(when_Stream_l1279) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 2'b01);
        if(when_Stream_l1314) begin
          logic_ptr_push <= 2'b00;
        end
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 2'b01);
        if(when_Stream_l1318) begin
          logic_ptr_pop <= 2'b00;
        end
      end
      if(io_flush) begin
        logic_ptr_push <= 2'b00;
        logic_ptr_pop <= 2'b00;
      end
      logic_ptr_notPow2_counter <= (_zz_logic_ptr_notPow2_counter - _zz_logic_ptr_notPow2_counter_3);
      if(io_flush) begin
        logic_ptr_notPow2_counter <= 2'b00;
      end
    end
  end


endmodule
